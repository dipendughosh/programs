TTLINV CKT - 74 SERIES TTL INVERTER

.MODEL D1 D(RS=40 TT=0.1NS CJO=0.9PF)
.MODEL QND NPN(BF=50 RB=70 RC=40 CCS=2PF TF=0.1NS TR=10NS
+ CJE=0.9PF CJC=1.5PF PC=0.85 VA=50)

VCC 13 0 5.0
VIN 1 0 PULSE(0 3.5 1NS 1NS 1NS 40NS)
RS 1 2 50
Q1 4 3 2 QND
RB1 13 3 4K
Q2 5 4 6 QND
RC2 13 5 1.4K
RE2 6 0 1K
Q3 7 5 8 QND
RC3 13 7 100
D1 8 9 D1
Q4 9 6 0 QND
Q5 11 10 9 QND
RB5 13 10 4K
D2 11 12 D1
D3 12 0 D1


.TRAN 1NS 100NS
.PRINT TRAN V(1) V(5) V(9)
.END
