MECLIII CKT - MOTOROLA MECL III ECL GATE

.MODEL D1 D(RS=40 TT=0.1NS CJO=0.9PF)
.MODEL QND NPN(BF=50 RB=70 RC=40 CCS=2PF TF=0.1NS TR=10NS
+ CJE=0.9PF CJC=1.5PF PC=0.85 VA=50)

VEE 22 0 -6.0
VIN 1 0 PULSE(-0.8 -1.8 0.2NS 0.2NS 0.2NS 10NS)

RS 1 2 50
Q1 4 2 6 QND
Q2 4 3 6 QND
Q3 5 7 6 QND
Q4 0 8 7 QND
D1 8 9 D1
D2 9 10 D1
RP1 3 22 50K
RC1 0 4 100
RC2 0 5 112
RE 6 22 380
R1 7 22 2K
R2 0 8 350
R3 10 22 1958
Q5 0 5 11 QND
Q6 0 4 12 QND
RP2 11 22 560
RP3 12 22 560
Q7 13 12 15 QND
Q8 14 16 15 QND
RE2 15 22 380
RC3 0 13 100
RC4 0 14 112
Q9 0 17 16 QND
R4 16 22 2K
R5 0 17 350
D3 17 18 D1
D4 18 19 D1
R6 19 22 1958
Q10 0 14 20 QND
Q11 0 13 21 QND
RP4 20 22 560
RP5 21 22 560

.TRAN 0.1NS 20NS
.PRINT TRAN V(1) V(12) V(21)
.END
