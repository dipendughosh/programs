1*******020689 ********  SPICE 2G.6    3/15/83 ********18:18:45*****

0* ECL CKT - EMITTER COUPLED LOGIC INVERTER                                      

0****     INPUT LISTING                    TEMPERATURE =   27.000 DEG C

0***********************************************************************




 Q1 3 2 4 0 QSTD 
 Q2 5 6 4 0 QSTD 
 Q3 8 5 7 0 QSTD 
 Q4 8 5 7 0 QSTD 
 RIN 1 2 50      
 RC1 8 3 120     
 RC2 8 5 135     
 RE 4 0 340      
 RTH1 7 0 125    
 RTH2 7 0 85     
 CLOAD 7 0 5P    
         
 *.MODEL QSTD NPN BF=80 RB=100 TF=0.3N TR=6N CJE=3P CJC=2P VAF=50
 *+ RBM=50 IRB=1.0E-3    
         
 .MODEL QSTD NPN IS=2E-16 BF=50 BR=0.1 RB=100 RC=10 TF=0.12N     
 +  TR=5N CJE=0.4P VJE=0.8 MJE=0.4 CJC=0.5P VJC=0.8 MJC=0.333    
 +  CJS=3P VAF=50 RBM=50 IRB=1.0E-4      
         
 VIN 1 0 PULSE(4.0 3.2 1NS 1NS 8NS 20NS) 
 VCC 8 0 5.0     
 VREF 6 0 3.6    
         
 .OPTIONS ABSTOL=1E-12 RELTOL=1E-5       
 .TRAN 0.25NS 50NS       
 .PRINT TRAN V(1,0) I(VIN) V(3,0) V(5,0) 
 .END    
1****************020689 ************************  SPICE 2G.6    3/15/83 ************************18:18:45****************

0* ECL CKT - EMITTER COUPLED LOGIC INVERTER                                      
0****                 BJT MODEL PARAMETERS                                 TEMPERATURE =   27.000 DEG C

0*************************************************************************************************************************




             QSTD    
0TYPE        NPN   
0IS        2.00d-16
0BF          50.000
0NF           1.000
0VAF       5.00d+01
0BR           0.100
0NR           1.000
0RB         100.000
0IRB       1.00d-04
0RBM         50.000
0RC          10.000
0CJE       4.00d-13
0VJE          0.800
0MJE          0.400
0TF        1.20d-10
0CJC       5.00d-13
0VJC          0.800
0MJC          0.333
0TR        5.00d-09
0CJS       3.00d-12
1****************020689 ************************  SPICE 2G.6    3/15/83 ************************18:18:45****************

0* ECL CKT - EMITTER COUPLED LOGIC INVERTER                                      
0****                 INITIAL TRANSIENT SOLUTION                           TEMPERATURE =   27.000 DEG C

0*************************************************************************************************************************


  NODE   VOLTAGE     NODE   VOLTAGE     NODE   VOLTAGE     NODE   VOLTAGE     NODE   VOLTAGE     NODE   VOLTAGE     NODE   VOLTAGE


 (  1)    4.0000    (  2)    3.9908    (  3)    3.9051    (  4)    3.1644    (  5)    4.7955    (  6)    3.6000    (  7)    3.8983

 (  8)    5.0000    




     VOLTAGE SOURCE CURRENTS

     NAME       CURRENT


     VIN      -1.831d-04

     VCC      -8.617d-02

     VREF     -7.069d-11


     TOTAL POWER DISSIPATION   4.32d-01  WATTS
1****************020689 ************************  SPICE 2G.6    3/15/83 ************************18:18:45****************

0* ECL CKT - EMITTER COUPLED LOGIC INVERTER                                      
0****                 OPERATING POINT INFORMATION                          TEMPERATURE =   27.000 DEG C

0*************************************************************************************************************************


0
0**** BIPOLAR JUNCTION TRANSISTORS


0            Q1        Q2        Q3        Q4      
0MODEL     QSTD      QSTD      QSTD      QSTD    
 IB        1.83e-04  7.07e-11  7.57e-04  7.57e-04
 IC        9.12e-03  4.24e-09  3.78e-02  3.78e-02
 VBE          0.826     0.436     0.897     0.897
 VBC          0.086    -1.196    -0.204    -0.204
 VCE          0.741     1.631     1.102     1.102
 BETADC      49.836    60.044    49.874    49.874
1****************020689 ************************  SPICE 2G.6    3/15/83 ************************18:18:45****************

0* ECL CKT - EMITTER COUPLED LOGIC INVERTER                                      
0****                 TRANSIENT ANALYSIS                                   TEMPERATURE =   27.000 DEG C

0*************************************************************************************************************************



     TIME       V(1)        I(VIN)      V(3)        V(5)        
X
 
  0.000e+00     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  2.500e-10     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  5.000e-10     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  7.500e-10     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  1.000e-09     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  1.250e-09     3.800e+00   4.816e-04   3.900e+00   4.794e+00
  1.500e-09     3.600e+00   6.371e-04   3.922e+00   4.793e+00
  1.750e-09     3.400e+00   1.241e-03   3.991e+00   4.773e+00
  2.000e-09     3.200e+00   2.069e-03   4.142e+00   4.698e+00
  2.250e-09     3.200e+00   1.711e-03   4.388e+00   4.559e+00
  2.500e-09     3.200e+00   1.049e-03   4.630e+00   4.388e+00
  2.750e-09     3.200e+00   4.200e-04   4.784e+00   4.236e+00
  3.000e-09     3.200e+00   1.774e-04   4.876e+00   4.118e+00
  3.250e-09     3.200e+00   8.997e-05   4.930e+00   4.029e+00
  3.500e-09     3.200e+00   5.204e-05   4.960e+00   3.964e+00
  3.750e-09     3.200e+00   3.041e-05   4.978e+00   3.915e+00
  4.000e-09     3.200e+00   1.826e-05   4.987e+00   3.878e+00
  4.250e-09     3.200e+00   1.088e-05   4.993e+00   3.851e+00
  4.500e-09     3.200e+00   6.523e-06   4.996e+00   3.830e+00
  4.750e-09     3.200e+00   4.069e-06   4.998e+00   3.815e+00
  5.000e-09     3.200e+00   2.563e-06   4.999e+00   3.804e+00
  5.250e-09     3.200e+00   1.638e-06   4.999e+00   3.795e+00
  5.500e-09     3.200e+00   1.068e-06   5.000e+00   3.789e+00
  5.750e-09     3.200e+00   7.124e-07   5.000e+00   3.784e+00
  6.000e-09     3.200e+00   4.857e-07   5.000e+00   3.781e+00
  6.250e-09     3.200e+00   3.371e-07   5.000e+00   3.778e+00
  6.500e-09     3.200e+00   2.365e-07   5.000e+00   3.776e+00
  6.750e-09     3.200e+00   1.662e-07   5.000e+00   3.774e+00
  7.000e-09     3.200e+00   1.196e-07   5.000e+00   3.773e+00
  7.250e-09     3.200e+00   8.810e-08   5.000e+00   3.772e+00
  7.500e-09     3.200e+00   6.288e-08   5.000e+00   3.772e+00
  7.750e-09     3.200e+00   4.720e-08   5.000e+00   3.771e+00
  8.000e-09     3.200e+00   3.421e-08   5.000e+00   3.771e+00
  8.250e-09     3.200e+00   2.579e-08   5.000e+00   3.771e+00
  8.500e-09     3.200e+00   1.846e-08   5.000e+00   3.770e+00
  8.750e-09     3.200e+00   1.427e-08   5.000e+00   3.770e+00
  9.000e-09     3.200e+00   1.008e-08   5.000e+00   3.770e+00
  9.250e-09     3.200e+00   7.689e-09   5.000e+00   3.770e+00
  9.500e-09     3.200e+00   5.861e-09   5.000e+00   3.770e+00
  9.750e-09     3.200e+00   4.034e-09   5.000e+00   3.770e+00
  1.000e-08     3.200e+00   3.049e-09   5.000e+00   3.770e+00
  1.025e-08     3.200e+00   2.387e-09   5.000e+00   3.770e+00
  1.050e-08     3.200e+00   1.724e-09   5.000e+00   3.770e+00
  1.075e-08     3.200e+00   1.062e-09   5.000e+00   3.770e+00
  1.100e-08     3.200e+00   8.249e-10   5.000e+00   3.770e+00
  1.125e-08     3.200e+00   6.405e-10   5.000e+00   3.770e+00
  1.150e-08     3.200e+00   4.560e-10   5.000e+00   3.770e+00
  1.175e-08     3.200e+00   2.715e-10   5.000e+00   3.770e+00
  1.200e-08     3.200e+00   2.045e-10   5.000e+00   3.770e+00
  1.225e-08     3.200e+00   1.521e-10   5.000e+00   3.770e+00
  1.250e-08     3.200e+00   9.968e-11   5.000e+00   3.770e+00
  1.275e-08     3.200e+00   4.728e-11   5.000e+00   3.770e+00
  1.300e-08     3.200e+00   3.063e-11   5.000e+00   3.770e+00
  1.325e-08     3.200e+00   1.842e-11   5.000e+00   3.770e+00
  1.350e-08     3.200e+00   6.222e-12   5.000e+00   3.770e+00
  1.375e-08     3.200e+00  -5.981e-12   5.000e+00   3.770e+00
  1.400e-08     3.200e+00  -1.180e-11   5.000e+00   3.770e+00
  1.425e-08     3.200e+00  -1.683e-11   5.000e+00   3.770e+00
  1.450e-08     3.200e+00  -2.186e-11   5.000e+00   3.770e+00
  1.475e-08     3.200e+00  -2.689e-11   5.000e+00   3.770e+00
  1.500e-08     3.200e+00   1.094e-12   5.000e+00   3.770e+00
  1.525e-08     3.200e+00   3.320e-11   5.000e+00   3.770e+00
  1.550e-08     3.200e+00   6.530e-11   5.000e+00   3.770e+00
  1.575e-08     3.200e+00   9.740e-11   5.000e+00   3.770e+00
  1.600e-08     3.200e+00   3.504e-12   5.000e+00   3.770e+00
  1.625e-08     3.200e+00  -1.061e-10   5.000e+00   3.770e+00
  1.650e-08     3.200e+00  -2.157e-10   5.000e+00   3.770e+00
  1.675e-08     3.200e+00  -3.253e-10   5.000e+00   3.770e+00
  1.700e-08     3.200e+00  -1.927e-10   5.000e+00   3.770e+00
  1.725e-08     3.200e+00  -2.985e-11   5.000e+00   3.770e+00
  1.750e-08     3.200e+00   1.330e-10   5.000e+00   3.770e+00
  1.775e-08     3.200e+00   2.958e-10   5.000e+00   3.770e+00
  1.800e-08     3.200e+00   1.410e-10   5.000e+00   3.770e+00
  1.825e-08     3.200e+00  -5.344e-11   5.000e+00   3.770e+00
  1.850e-08     3.200e+00  -2.479e-10   5.000e+00   3.770e+00
  1.875e-08     3.200e+00  -4.423e-10   5.000e+00   3.770e+00
  1.900e-08     3.200e+00  -2.396e-10   5.000e+00   3.770e+00
  1.925e-08     3.200e+00   1.267e-11   5.000e+00   3.770e+00
  1.950e-08     3.200e+00   2.649e-10   5.000e+00   3.770e+00
  1.975e-08     3.200e+00   5.172e-10   5.000e+00   3.770e+00
  2.000e-08     3.200e+00   2.922e-10   5.000e+00   3.770e+00
  2.025e-08     3.200e+00   7.766e-12   5.000e+00   3.770e+00
  2.050e-08     3.200e+00  -2.767e-10   5.000e+00   3.770e+00
  2.075e-08     3.200e+00  -5.612e-10   5.000e+00   3.770e+00
  2.100e-08     3.200e+00  -3.637e-10   5.000e+00   3.770e+00
  2.125e-08     3.200e+00  -1.061e-10   5.000e+00   3.770e+00
  2.150e-08     3.200e+00   1.515e-10   5.000e+00   3.770e+00
  2.175e-08     3.200e+00   4.090e-10   5.000e+00   3.770e+00
  2.200e-08     3.200e+00  -8.219e-10   5.000e+00   3.770e+00
  2.225e-08     3.225e+00  -7.194e-05   5.001e+00   3.770e+00
  2.250e-08     3.250e+00  -8.623e-05   5.002e+00   3.771e+00
  2.275e-08     3.275e+00  -8.966e-05   5.003e+00   3.773e+00
  2.300e-08     3.300e+00  -9.133e-05   5.003e+00   3.774e+00
  2.325e-08     3.325e+00  -9.293e-05   5.004e+00   3.774e+00
  2.350e-08     3.350e+00  -9.453e-05   5.004e+00   3.775e+00
  2.375e-08     3.375e+00  -9.634e-05   5.004e+00   3.776e+00
  2.400e-08     3.400e+00  -9.853e-05   5.004e+00   3.776e+00
  2.425e-08     3.425e+00  -1.016e-04   5.004e+00   3.777e+00
  2.450e-08     3.450e+00  -1.066e-04   5.003e+00   3.778e+00
  2.475e-08     3.475e+00  -1.160e-04   5.001e+00   3.779e+00
  2.500e-08     3.500e+00  -1.333e-04   4.998e+00   3.781e+00
  2.525e-08     3.525e+00  -1.629e-04   4.992e+00   3.785e+00
  2.550e-08     3.550e+00  -2.042e-04   4.980e+00   3.792e+00
  2.575e-08     3.575e+00  -2.573e-04   4.961e+00   3.804e+00
  2.600e-08     3.600e+00  -3.190e-04   4.934e+00   3.823e+00
  2.625e-08     3.625e+00  -3.879e-04   4.897e+00   3.849e+00
  2.650e-08     3.650e+00  -4.614e-04   4.849e+00   3.884e+00
  2.675e-08     3.675e+00  -5.371e-04   4.790e+00   3.929e+00
  2.700e-08     3.700e+00  -6.133e-04   4.721e+00   3.982e+00
  2.725e-08     3.725e+00  -6.855e-04   4.638e+00   4.050e+00
  2.750e-08     3.750e+00  -7.527e-04   4.549e+00   4.124e+00
  2.775e-08     3.775e+00  -8.075e-04   4.450e+00   4.208e+00
  2.800e-08     3.800e+00  -8.375e-04   4.345e+00   4.299e+00
  2.825e-08     3.825e+00  -8.046e-04   4.238e+00   4.395e+00
  2.850e-08     3.850e+00  -6.261e-04   4.141e+00   4.485e+00
  2.875e-08     3.875e+00  -4.218e-04   4.067e+00   4.559e+00
  2.900e-08     3.900e+00  -3.442e-04   4.017e+00   4.617e+00
  2.925e-08     3.925e+00  -3.190e-04   3.985e+00   4.661e+00
  2.950e-08     3.950e+00  -3.067e-04   3.963e+00   4.694e+00
  2.975e-08     3.975e+00  -2.998e-04   3.947e+00   4.719e+00
  3.000e-08     4.000e+00  -2.964e-04   3.935e+00   4.738e+00
  3.025e-08     4.000e+00  -2.123e-04   3.923e+00   4.752e+00
  3.050e-08     4.000e+00  -1.961e-04   3.916e+00   4.763e+00
  3.075e-08     4.000e+00  -1.912e-04   3.911e+00   4.771e+00
  3.100e-08     4.000e+00  -1.883e-04   3.909e+00   4.777e+00
  3.125e-08     4.000e+00  -1.863e-04   3.907e+00   4.781e+00
  3.150e-08     4.000e+00  -1.850e-04   3.906e+00   4.785e+00
  3.175e-08     4.000e+00  -1.842e-04   3.906e+00   4.788e+00
  3.200e-08     4.000e+00  -1.837e-04   3.906e+00   4.790e+00
  3.225e-08     4.000e+00  -1.834e-04   3.905e+00   4.791e+00
  3.250e-08     4.000e+00  -1.833e-04   3.905e+00   4.792e+00
  3.275e-08     4.000e+00  -1.832e-04   3.905e+00   4.793e+00
  3.300e-08     4.000e+00  -1.831e-04   3.905e+00   4.794e+00
  3.325e-08     4.000e+00  -1.831e-04   3.905e+00   4.794e+00
  3.350e-08     4.000e+00  -1.831e-04   3.905e+00   4.794e+00
  3.375e-08     4.000e+00  -1.831e-04   3.905e+00   4.795e+00
  3.400e-08     4.000e+00  -1.831e-04   3.905e+00   4.795e+00
  3.425e-08     4.000e+00  -1.831e-04   3.905e+00   4.795e+00
  3.450e-08     4.000e+00  -1.831e-04   3.905e+00   4.795e+00
  3.475e-08     4.000e+00  -1.831e-04   3.905e+00   4.795e+00
  3.500e-08     4.000e+00  -1.831e-04   3.905e+00   4.795e+00
  3.525e-08     4.000e+00  -1.831e-04   3.905e+00   4.795e+00
  3.550e-08     4.000e+00  -1.831e-04   3.905e+00   4.795e+00
  3.575e-08     4.000e+00  -1.831e-04   3.905e+00   4.795e+00
  3.600e-08     4.000e+00  -1.831e-04   3.905e+00   4.795e+00
  3.625e-08     4.000e+00  -1.831e-04   3.905e+00   4.795e+00
  3.650e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  3.675e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  3.700e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  3.725e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  3.750e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  3.775e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  3.800e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  3.825e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  3.850e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  3.875e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  3.900e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  3.925e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  3.950e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  3.975e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.000e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.025e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.050e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.075e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.100e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.125e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.150e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.175e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.200e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.225e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.250e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.275e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.300e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.325e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.350e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.375e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.400e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.425e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.450e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.475e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.500e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.525e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.550e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.575e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.600e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.625e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.650e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.675e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.700e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.725e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.750e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.775e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.800e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.825e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.850e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.875e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.900e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.925e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.950e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  4.975e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
  5.000e-08     4.000e+00  -1.831e-04   3.905e+00   4.796e+00
Y
0
         JOB CONCLUDED
0         TOTAL JOB TIME           16.17
