magic
tech hpcmos40
timestamp 588531989
<< ndiffusion >>
rect -21 8 79 17
rect 83 8 283 17
rect 290 8 690 17
rect -21 3 79 4
rect 83 3 283 4
rect 290 3 690 4
<< pdiffusion >>
rect -21 -32 79 -31
rect 83 -32 283 -31
rect 290 -32 690 -31
rect -21 -45 79 -36
rect 83 -45 283 -36
rect 290 -45 690 -36
<< polysilicon >>
rect -30 4 -21 8
rect 79 4 83 8
rect 283 4 290 8
rect 690 4 694 8
rect -30 3 -22 4
rect -30 -32 -22 -31
rect -30 -36 -21 -32
rect 79 -36 83 -32
rect 283 -36 290 -32
rect 690 -36 695 -32
<< metal1 >>
rect -22 -5 -21 3
rect 79 -5 83 3
rect 283 -5 290 3
rect -22 -31 -21 -23
rect 79 -31 83 -23
rect 283 -31 290 -23
<< polycontact >>
rect -30 -5 -22 3
rect -30 -31 -22 -23
<< ndcontact >>
rect -21 -5 79 3
rect 83 -5 283 3
rect 290 -5 690 3
<< pdcontact >>
rect -21 -31 79 -23
rect 83 -31 283 -23
rect 290 -31 690 -23
<< ntransistor >>
rect -21 4 79 8
rect 83 4 283 8
rect 290 4 690 8
<< ptransistor >>
rect -21 -36 79 -32
rect 83 -36 283 -32
rect 290 -36 690 -32
<< labels >>
rlabel ndiffusion -17 15 -17 15 5 drain1
rlabel pdiffusion -16 -44 -16 -44 1 drain4
rlabel ndiffusion 91 15 91 15 5 drain2
rlabel pdiffusion 91 -44 91 -44 1 drain5
rlabel metal1 288 -1 288 -1 1 GND
rlabel ndiffusion 309 14 309 14 5 drain3
rlabel pdiffusion 310 -44 310 -44 1 drain6
rlabel metal1 286 -27 286 -27 1 Vdd
<< end >>
