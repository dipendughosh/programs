SCHMITT CKT - ECL COMPATIBLE SCHMITT TRIGGER

.MODEL QSTD NPN
+ is=1E-16 BF=50 BR=0.1 RB=50 RC=10 TF=0.12N
+   TR=5NS CJE=0.4P PE=0.8 ME=0.4 CJC=0.5P PC=0.8 MC=0.333
+   CCS=1p VA=50

VIN 1 0 PULSE(-1.6 -1.2 10ns 400ns 400ns 100ns 1000ns )
VEE 8 0 -5.0
RIN 1 2 50
RC1 0 3 50
R1 3 5 185
R2 5 8 760
RC2 0 6 100
RE 4 8 260
RTH1 7 8 125
RTH2 7 0 85
CLOAD 7 0 5P
Q1 3 2 4 QSTD OFF
Q2 6 5 4 QSTD
Q3 8 6 7 QSTD
Q4 8 6 7 QSTD


.print tran v(1) v(3) v(5) v(6)
.tran 10ns 1000ns
.option acct limpts=100000 numdgt=6
.end
 
