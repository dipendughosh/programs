RC CKT - SPLIT TIME-CONSTANT RC CIRCUIT
VIN 1 0 PULSE(0 1 0.1MS 0.1MS)
R1 1 2 1K
C1 2 0 1PF
R2 2 3 1K
C2 3 0 1UF
.TRAN 0.1MS 10MS
.PRINT TRAN V(1) V(2) V(3)
.END

