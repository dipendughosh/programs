sig.sp SPICE FILE
.model nenh nmos
+ level = 2
+    vto = 0.779   kp = 3.52e-05   gamma = 1.04
+    phi = 0.6
+ 
+    cgso = 5.2e-10   cgdo = 5.2e-10
+    rsh = 25   cj = 0.00042
+    mj = 0.5   cjsw = 9e-10   mjsw = 0.33
+    tox = 5e-08   nsub = 1e+16
+    nss = 0   nfs = 1.306e+11   tpg = 1
+    xj = 3.85e-08   ld = 1e-07   uo = 400
+    ucrit = 999000   uexp = 0.001001
+    vmax = 32585.3   neff = 0.01001
+ 
+    delta = 1.33
.model penh pmos
+ level = 2
+    vto = -0.988   kp = 1.206e-05   gamma = 0.619
+    phi = 0.6
+ 
+    cgso = 4e-10   cgdo = 4e-10
+    rsh = 95   cj = 0.00032
+    mj = 0.5   cjsw = 5.5e-10   mjsw = 0.33
+    tox = 5e-08   nsub = 8.158e+14
+    nss = 0   nfs = 5.55e+09   tpg = -1
+    xj = 1.46e-07   ld = 2.52e-07   uo = 150
+    ucrit = 54941   uexp = 0.17
+    vmax = 100000   neff = 0.01001
+ 
+    delta = 1.129
mm2 3 4 1 1 penh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm3 3 4 0 0 nenh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm4 5 6 1 1 penh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm5 5 6 0 0 nenh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm6 7 8 1 1 penh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm7 7 8 0 0 nenh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm8 9 10 1 1 penh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm9 9 10 0 0 nenh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm12 11 12 1 1 penh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm13 11 12 0 0 nenh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm14 13 14 1 1 penh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm15 13 14 0 0 nenh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm16 15 16 1 1 penh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm17 15 16 0 0 nenh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm18 17 18 1 1 penh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm19 17 18 0 0 nenh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm20 19 20 1 1 penh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm21 19 20 0 0 nenh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm22 21 22 1 1 penh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
mm23 21 22 0 0 nenh l=3e-06 w=7e-06 as=5.6e-11 ad=5.6e-11 
+ ps=3e-05 pd=3e-05 nrd=1e-30 nrs=1e-30
rR1 23 0 1000
rR2 24 0 1000
Vvdd 0 0 5
Vf0 4 0 pwl (0 5 1.999e-06 5 2e-06 0 1.5999e-05 0 1.6e-05 5 
+ 1.7999e-05 5 1.8e-05 0 1.9999e-05 0 2e-05 5 2.1999e-05 5 
+ 2.3999e-05 0 3.9998e-05 0 5.5998e-05 5 7.3997e-05 5 9.1997e-05 0 
+ )
Vf1 6 0 pwl (0 0 1.999e-06 0 2e-06 5 3.999e-06 5 4e-06 0 
+ 1.7999e-05 0 1.8e-05 5 1.9999e-05 5 2e-05 0 2.1999e-05 0 
+ 2.3999e-05 5 2.7998e-05 5 3.1998e-05 0 4.9997e-05 0 6.7997e-05 5 
+ 8.7996e-05 5 )
Vf2 8 0 pwl (0 0 4e-06 0 4.001e-06 5 6e-06 5 6.001e-06 0 
+ 2e-05 0 2.4e-05 0 2.8001e-05 5 3.4001e-05 5 4.0002e-05 0 
+ 6.0002e-05 0 6.4002e-05 0 6.8003e-05 5 7.4003e-05 5 8.0004e-05 0 
+ )
Vf3 10 0 pwl (0 0 1e-05 0 1.0001e-05 5 1.2e-05 5 1.2001e-05 0 
+ 2e-05 0 3e-05 0 4.0001e-05 5 5.2001e-05 5 6.4002e-05 0 
+ 8.4002e-05 0 )
Vcltc 22 0 pwl (0 0 2e-06 5 4e-06 5 8e-06 0 1e-05 5 
+ 1.4e-05 5 2.2e-05 0 2.4e-05 5 2.8e-05 5 3.6e-05 0 
+ 3.8e-05 5 4.2e-05 5 5e-05 0 5.2e-05 5 5.6e-05 5 
+ 6.4e-05 0 6.6e-05 5 7e-05 5 7.8e-05 0 8e-05 5 
+ )
Vcltx 12 0 pwl (0 0 2.49e-07 0 2.5e-07 5 4.99e-07 5 5e-07 0 
+ 7.49e-07 0 9.99e-07 5 1.498e-06 5 1.998e-06 0 2.247e-06 0 
+ 2.497e-06 5 2.996e-06 5 3.496e-06 0 3.745e-06 0 3.995e-06 5 
+ 4.494e-06 5 4.994e-06 0 5.243e-06 0 5.493e-06 5 5.992e-06 5 
+ 6.492e-06 0 6.741e-06 0 6.991e-06 5 7.49e-06 5 7.99e-06 0 
+ 8.239e-06 0 8.489e-06 5 8.988e-06 5 9.488e-06 0 9.737e-06 0 
+ 9.987e-06 5 1.0486e-05 5 1.0986e-05 0 1.1235e-05 0 1.1485e-05 5 
+ 1.1984e-05 5 1.2484e-05 0 1.2733e-05 0 1.2983e-05 5 1.3482e-05 5 
+ 1.3982e-05 0 1.4231e-05 0 1.4481e-05 5 1.498e-05 5 1.548e-05 0 
+ 1.5729e-05 0 1.5979e-05 5 1.6478e-05 5 1.6978e-05 0 1.7227e-05 0 
+ 1.7477e-05 5 1.7976e-05 5 1.8476e-05 0 1.8725e-05 0 1.8975e-05 5 
+ 1.9474e-05 5 1.9974e-05 0 2.0223e-05 0 2.0473e-05 5 2.0972e-05 5 
+ 2.1472e-05 0 2.1721e-05 0 2.1971e-05 5 2.247e-05 5 2.297e-05 0 
+ 2.3219e-05 0 2.3469e-05 5 2.3968e-05 5 2.4468e-05 0 2.4717e-05 0 
+ 2.4967e-05 5 2.5466e-05 5 2.5966e-05 0 2.6215e-05 0 2.6465e-05 5 
+ 2.6964e-05 5 2.7464e-05 0 2.7713e-05 0 2.7963e-05 5 2.8462e-05 5 
+ 2.8962e-05 0 2.9211e-05 0 2.9461e-05 5 2.996e-05 5 3.046e-05 0 
+ 3.0709e-05 0 3.0959e-05 5 3.1458e-05 5 3.1958e-05 0 3.2207e-05 0 
+ 3.2457e-05 5 3.2956e-05 5 3.3456e-05 0 3.3705e-05 0 3.3955e-05 5 
+ 3.4454e-05 5 3.4954e-05 0 3.5203e-05 0 3.5453e-05 5 3.5952e-05 5 
+ 3.6452e-05 0 3.6701e-05 0 3.6951e-05 5 3.745e-05 5 3.795e-05 0 
+ 3.8199e-05 0 3.8449e-05 5 3.8948e-05 5 3.9448e-05 0 3.9697e-05 0 
+ 3.9947e-05 5 4.0446e-05 5 4.0946e-05 0 4.1195e-05 0 4.1445e-05 5 
+ 4.1944e-05 5 4.2444e-05 0 4.2693e-05 0 4.2943e-05 5 4.3442e-05 5 
+ 4.3942e-05 0 4.4191e-05 0 4.4441e-05 5 4.494e-05 5 4.544e-05 0 
+ 4.5689e-05 0 4.5939e-05 5 4.6438e-05 5 4.6938e-05 0 4.7187e-05 0 
+ 4.7437e-05 5 4.7936e-05 5 4.8436e-05 0 4.8685e-05 0 4.8935e-05 5 
+ 4.9434e-05 5 4.9934e-05 0 5.0183e-05 0 5.0433e-05 5 5.0932e-05 5 
+ 5.1432e-05 0 5.1681e-05 0 5.1931e-05 5 5.243e-05 5 5.293e-05 0 
+ 5.3179e-05 0 5.3429e-05 5 5.3928e-05 5 5.4428e-05 0 5.4677e-05 0 
+ 5.4927e-05 5 5.5426e-05 5 5.5926e-05 0 5.6175e-05 0 5.6425e-05 5 
+ 5.6924e-05 5 5.7424e-05 0 5.7673e-05 0 5.7923e-05 5 5.8422e-05 5 
+ 5.8922e-05 0 5.9171e-05 0 5.9421e-05 5 5.992e-05 5 6.042e-05 0 
+ 6.0669e-05 0 6.0919e-05 5 6.1418e-05 5 6.1918e-05 0 6.2167e-05 0 
+ 6.2417e-05 5 6.2916e-05 5 6.3416e-05 0 6.3665e-05 0 6.3915e-05 5 
+ 6.4414e-05 5 6.4914e-05 0 6.5163e-05 0 6.5413e-05 5 6.5912e-05 5 
+ 6.6412e-05 0 6.6661e-05 0 6.6911e-05 5 6.741e-05 5 6.791e-05 0 
+ 6.8159e-05 0 6.8409e-05 5 6.8908e-05 5 6.9408e-05 0 6.9657e-05 0 
+ 6.9907e-05 5 7.0406e-05 5 7.0906e-05 0 7.1155e-05 0 7.1405e-05 5 
+ 7.1904e-05 5 7.2404e-05 0 7.2653e-05 0 7.2903e-05 5 7.3402e-05 5 
+ 7.3902e-05 0 7.4151e-05 0 7.4401e-05 5 7.49e-05 5 7.54e-05 0 
+ 7.5649e-05 0 7.5899e-05 5 7.6398e-05 5 7.6898e-05 0 7.7147e-05 0 
+ 7.7397e-05 5 7.7896e-05 5 7.8396e-05 0 7.8645e-05 0 7.8895e-05 5 
+ 7.9394e-05 5 7.9894e-05 0 8.0143e-05 0 )
Vclty 14 0 pwl (0 0 4.99e-07 0 5e-07 5 9.99e-07 5 1e-06 0 
+ 1.499e-06 0 1.999e-06 5 2.998e-06 5 3.998e-06 0 4.497e-06 0 
+ 4.997e-06 5 5.996e-06 5 6.996e-06 0 7.495e-06 0 7.995e-06 5 
+ 8.994e-06 5 9.994e-06 0 1.0493e-05 0 1.0993e-05 5 1.1992e-05 5 
+ 1.2992e-05 0 1.3491e-05 0 1.3991e-05 5 1.499e-05 5 1.599e-05 0 
+ 1.6489e-05 0 1.6989e-05 5 1.7988e-05 5 1.8988e-05 0 1.9487e-05 0 
+ 1.9987e-05 5 2.0986e-05 5 2.1986e-05 0 2.2485e-05 0 2.2985e-05 5 
+ 2.3984e-05 5 2.4984e-05 0 2.5483e-05 0 2.5983e-05 5 2.6982e-05 5 
+ 2.7982e-05 0 2.8481e-05 0 2.8981e-05 5 2.998e-05 5 3.098e-05 0 
+ 3.1479e-05 0 3.1979e-05 5 3.2978e-05 5 3.3978e-05 0 3.4477e-05 0 
+ 3.4977e-05 5 3.5976e-05 5 3.6976e-05 0 3.7475e-05 0 3.7975e-05 5 
+ 3.8974e-05 5 3.9974e-05 0 4.0473e-05 0 4.0973e-05 5 4.1972e-05 5 
+ 4.2972e-05 0 4.3471e-05 0 4.3971e-05 5 4.497e-05 5 4.597e-05 0 
+ 4.6469e-05 0 4.6969e-05 5 4.7968e-05 5 4.8968e-05 0 4.9467e-05 0 
+ 4.9967e-05 5 5.0966e-05 5 5.1966e-05 0 5.2465e-05 0 5.2965e-05 5 
+ 5.3964e-05 5 5.4964e-05 0 5.5463e-05 0 5.5963e-05 5 5.6962e-05 5 
+ 5.7962e-05 0 5.8461e-05 0 5.8961e-05 5 5.996e-05 5 6.096e-05 0 
+ 6.1459e-05 0 6.1959e-05 5 6.2958e-05 5 6.3958e-05 0 6.4457e-05 0 
+ 6.4957e-05 5 6.5956e-05 5 6.6956e-05 0 6.7455e-05 0 6.7955e-05 5 
+ 6.8954e-05 5 6.9954e-05 0 7.0453e-05 0 7.0953e-05 5 7.1952e-05 5 
+ 7.2952e-05 0 7.3451e-05 0 7.3951e-05 5 7.495e-05 5 7.595e-05 0 
+ 7.6449e-05 0 7.6949e-05 5 7.7948e-05 5 7.8948e-05 0 7.9447e-05 0 
+ 7.9947e-05 5 8.0946e-05 5 )
Icltz 16 0 pwl (0 0 9.99e-07 0 1e-06 5e-06 1.999e-06 5e-06 2e-06 0 
+ 2.999e-06 0 3.999e-06 5e-06 5.998e-06 5e-06 7.998e-06 0 8.997e-06 0 
+ 9.997e-06 5e-06 1.1996e-05 5e-06 1.3996e-05 0 1.4995e-05 0 1.5995e-05 5e-06 
+ 1.7994e-05 5e-06 1.9994e-05 0 2.0993e-05 0 2.1993e-05 5e-06 2.3992e-05 5e-06 
+ 2.5992e-05 0 2.6991e-05 0 2.7991e-05 5e-06 2.999e-05 5e-06 3.199e-05 0 
+ 3.2989e-05 0 3.3989e-05 5e-06 3.5988e-05 5e-06 3.7988e-05 0 3.8987e-05 0 
+ 3.9987e-05 5e-06 4.1986e-05 5e-06 4.3986e-05 0 4.4985e-05 0 4.5985e-05 5e-06 
+ 4.7984e-05 5e-06 4.9984e-05 0 5.0983e-05 0 5.1983e-05 5e-06 5.3982e-05 5e-06 
+ 5.5982e-05 0 5.6981e-05 0 5.7981e-05 5e-06 5.998e-05 5e-06 6.198e-05 0 
+ 6.2979e-05 0 6.3979e-05 5e-06 6.5978e-05 5e-06 6.7978e-05 0 6.8977e-05 0 
+ 6.9977e-05 5e-06 7.1976e-05 5e-06 7.3976e-05 0 7.4975e-05 0 7.5975e-05 5e-06 
+ 7.7974e-05 5e-06 7.9974e-05 0 8.0973e-05 0 )
Vgg 18 25 (0.5 2 1e+07 0 0 )
Icltb 20 0 (5e-07 2e-06 1e+07 0 0 )
.options reltol=1e-07 abstol=5e-10 chgtol=5e-15 numdgt = 4 limpts = 10000
.print TRAN v(18) v(20) v(22) 
.print TRAN v(4) v(6) v(8) v(10) v(12) v(14) v(16) 
.TRAN 1e-07 8e-05
.end
