TL FOR ADDRESS SIGNAL         
.SUBCKT TL 22 500  42       
R11 22 23 0.10588   
R12 24 25 0.10588   
R13 26 27 0.10588   
R14 28 29 0.10588   
R15 30 31 0.10588   
R16 32 33 0.10588   
R17 34 35 0.10588   
R18 36 37 0.10588   
R19 38 39 0.10588   
R20 40 41 0.10588   
L11 23 24 0.2497NH  
L12 25 26 0.2497NH  
L13 27 28 0.2497NH  
L14 29 30 0.2497NH  
L15 31 32 0.2497NH  
L16 33 34 0.2497NH  
L17 35 36 0.2497NH  
L18 37 38 0.2497NH  
L19 39 40 0.2497NH  
L20 41 42 0.2497NH  
C11 24 500 0.15604PF
C12 26 500 0.15604PF
C13 28 500 0.15604PF
C14 30 500 0.15604PF
C15 32 500 0.15604PF
C16 34 500 0.15604PF
C17 36 500 0.15604PF
C18 38 500 0.15604PF
C19 40 500 0.15604PF
C20 42 500 0.15604PF
.ENDS TL    
.SUBCKT SB 901 99 90
C901 901 99 0.4PF   
C90 90 99 0.4PF     
L901 901 90 0.1NH   
.ENDS SB    
X1 20 0 1120 TL     
X2 1120 0 1220 TL   
X3 1220 0 1320 TL   
X4 1320 0 1420 TL   
X5 1420 0 1520 TL   
X6 1520 0 1620 TL   
X7 1620 0 1720 TL   
X8 1720 0 203 TL    
X22 1120 0 1121 SB  
R220 1121 0 1000K   
C220 1121 0 2.5PF    
X25 1220 0 1221 SB  
R250 1221 0 1000K   
C250 1220 0 2.5PF    
X28 1320 0 1321 SB  
R280 1321 0 1000K   
C280 1321 0 2.5PF    
X31 1420 0 1421 SB  
R310 1421 0 1000K   
C310 1421 0 2.5PF    
X34 1520 0 1521 SB  
R340 1521 0 1000K   
C340 1521 0 2.5PF    
X37 1620 0 1621 SB  
R370 1621 0 1000K   
C370 1621 0 2.5PF    
X40 1720 0 1721 SB  
R400 1721 0 1000K   
C400 1721 0 2.5PF    
C201 201 0 0.4PF    
C20 20 0 0.4PF      
C203 203 0 0.4PF    
C204 204 0 0.4PF    
L201 201 20 0.1NH   
L203 203 204 0.1NH  
*   
** OUTPUT IMPEDANCE 
*   
CMODUL2 204 0 2.5PF 
*********************************************************** 
**************************************************************      
**	SECOND ROW       
*********************************************************** 
X21 50 0 1150 TL    
XR22 1150 0 1250 TL 
X23 1250 0 1350 TL  
X24 1350 0 1450 TL  
XR25 1450 0 1550 TL 
X26 1550 0 1650 TL  
X27 1650 0 1750 TL  
XR28 1750 0 213 TL  
X222 1150 0 1121 SB 
R2220 1121 0 1000K  
C2220 1121 0 2.5PF   
X225 1250 0 1251 SB 
R2250 1251 0 1000K  
C2250 1251 0 2.5PF   
X228 1350 0 1351 SB 
R2280 1351 0 1000K  
C2280 1351 0 2.5PF   
X231 1450 0 1451 SB 
R2310 1451 0 1000K  
C2310 1451 0 2.5PF   
X234 1550 0 1551 SB 
R2340 1551 0 1000K  
C2340 1551 0 2.5PF   
X237 1650 0 1651 SB 
R2370 1651 0 1000K  
C2370 1651 0 2.5PF   
X240 1750 0 1751 SB 
R2400 1751 0 1000K  
C2400 1751 0 2.5PF   
C2201 51 0 0.4PF    
CR220 50 0 0.4PF    
C2203 213 0 0.4PF   
C2204 214 0 0.4PF   
L2201 51 50 0.1NH   
L2203 213 214 0.1NH 
*   
** OUTPUT IMPEDANC2E
*   
C2MODUL22 214 0 2.5PF       
*********************************************************** 
**************************************************************      
***	THIRD ROW       
*********************************************************** 
XR31 80 0 1180 TL   
X32 1180 0 1280 TL  
X33 1280 0 1380 TL  
XR34 1380 0 1480 TL 
X35 1480 0 1580 TL  
X36 1580 0 1680 TL  
XR37 1680 0 1780 TL 
X38 1780 0 223 TL   
X322 1180 0 1181 SB 
R3220 1181 0 1000K  
C3220 1181 0 2.5PF   
X325 1280 0 1281 SB 
R3250 1281 0 1000K  
C3250 1281 0 2.5PF   
X328 1380 0 1381 SB 
R3280 1381 0 1000K  
C3280 1381 0 2.5PF   
X331 1480 0 1481 SB 
R3310 1481 0 1000K  
C3310 1481 0 2.5PF   
X334 1580 0 1581 SB 
R3340 1581 0 1000K  
C3340 1581 0 2.5PF   
X337 1680 0 1681 SB 
R3370 1681 0 1000K  
C3370 1681 0 2.5PF   
X340 1780 0 1781 SB 
R3400 1781 0 1000K  
C3400 1781 0 2.5PF   
C3201 1021 0 0.4PF  
C320 80 0 0.4PF     
C3203 223 0 0.4PF   
C3204 224 0 0.4PF   
L3201 1021 80 0.1NH 
L3203 223 224 0.1NH 
*   
** OUTPUT IMPEDANC3E
*   
C3MODUL32 224 0 2.5PF       
*********************************************************** 
**************************************************************      
***	4TH ROW 
*********************************************************** 
X41 1020 0 2120 TL  
X42 2120 0 2220 TL  
X43 2220 0 2320 TL  
X44 2320 0 2420 TL  
X45 2420 0 2520 TL  
X46 2520 0 2620 TL  
X47 2620 0 2720 TL  
X48 2720 0 233 TL   
X422 2120 0 2121 SB 
R4220 2121 0 1000K  
C4220 2121 0 2.5PF   
X425 2220 0 2221 SB 
R4250 2221 0 1000K  
C4250 2221 0 2.5PF   
X428 2320 0 2321 SB 
R4280 2321 0 1000K  
C4280 2321 0 2.5PF   
X431 2420 0 2421 SB 
R4310 2421 0 1000K  
C4310 2421 0 2.5PF   
X434 2520 0 2521 SB 
R4340 2521 0 1000K  
C4340 2521 0 2.5PF   
X437 2620 0 2621 SB 
R4370 2621 0 1000K  
C4370 2621 0 2.5PF   
X440 2720 0 2721 SB 
R4400 2721 0 1000K  
C4400 2721 0 2.5PF   
C4201 1021 0 0.4PF  
C420 1020 0 0.4PF   
C4203 233 0 0.4PF   
C4204 234 0 0.4PF   
L4201 1021 1020 0.1NH       
L4203 233 234 0.1NH 
*   
** OUTPUT IMPEDANC4E
*   
C4MODUL42 234 0 2.5PF       
*********************************************************** 
**************************************************************      
***	5TH ROW 
*********************************************************** 
X51 1050 0 2150 TL  
X52 2150 0 2250 TL  
X53 2250 0 2350 TL  
X54 2350 0 2450 TL  
X55 2450 0 2250 TL  
X56 2250 0 2650 TL  
X57 2650 0 2750 TL  
X58 2750 0 243 TL   
X522 2150 0 2151 SB 
R5220 2151 0 1000K  
C5220 2151 0 2.5PF   
X525 2250 0 2251 SB 
R5250 2251 0 1000K  
C5250 2251 0 2.5PF   
X528 2350 0 2351 SB 
R5280 2351 0 1000K  
C5280 2351 0 2.5PF   
X531 2450 0 2451 SB 
R5310 2451 0 1000K  
C5310 2451 0 2.5PF   
X534 2250 0 2551 SB 
R5340 2551 0 1000K  
C5340 2551 0 2.5PF   
X537 2650 0 2651 SB 
R5370 2651 0 1000K  
C5370 2651 0 2.5PF   
X540 2750 0 2751 SB 
R5400 2751 0 1000K  
C5400 2751 0 2.5PF   
C5201 1051 0 0.4PF  
C520 1050 0 0.4PF   
C5203 243 0 0.4PF   
C5204 244 0 0.4PF   
L5201 1051 1050 0.1NH       
L5203 243 244 0.1NH 
*   
** OUTPUT IMPEDANC5E
*   
C5MODUL52 244 0 2.5PF       
*********************************************************** 
**************************************************************      
***	6TH ROW 
*********************************************************** 
X61 1080 0 2180 TL  
X62 2180 0 2280 TL  
X63 2280 0 2380 TL  
X64 2380 0 2480 TL  
X65 2480 0 2580 TL  
X66 2580 0 2680 TL  
X67 2680 0 2780 TL  
X68 2780 0 253 TL   
X622 2180 0 2181 SB 
R6220 2181 0 1000K  
C6220 2181 0 2.5PF   
X625 2280 0 2281 SB 
R6250 2281 0 1000K  
C6250 2281 0 2.5PF   
X628 2380 0 2381 SB 
R6280 2381 0 1000K  
C6280 2381 0 2.5PF   
X631 2480 0 2481 SB 
R6310 2481 0 1000K  
C6310 2481 0 2.5PF   
X634 2580 0 2581 SB 
R6340 2581 0 1000K  
C6340 2581 0 2.5PF   
X637 2680 0 2681 SB 
R6370 2681 0 1000K  
C6370 2681 0 2.5PF   
X640 2780 0 2781 SB 
R6400 2781 0 1000K  
C6400 2781 0 2.5PF   
C6201 1081 0 0.4PF  
C620 1080 0 0.4PF   
C6203 253 0 0.4PF   
C6204 254 0 0.4PF   
L6201 1081 1080 0.1NH       
L6203 253 254 0.1NH 
*   
** OUTPUT IMPEDANC6E
*   
C6MODUL62 254 0 2.5PF       
*********************************************************** 
**************************************************************      
*** 7TH ROW 
*********************************************************** 
X71 2020 0 3120 TL  
X72 3120 0 3220 TL  
X73 3220 0 3320 TL  
X74 3320 0 3420 TL  
X75 3420 0 3520 TL  
X76 3520 0 3620 TL  
X77 3620 0 3720 TL  
X78 3720 0 263 TL   
X722 3120 0 3121 SB 
R7220 3121 0 1000K  
C7220 3121 0 2.5PF   
X725 3220 0 3221 SB 
R7250 3221 0 1000K  
C7250 3221 0 2.5PF   
X728 3320 0 3321 SB 
R7280 3321 0 1000K  
C7280 3321 0 2.5PF   
X731 3420 0 3421 SB 
R7310 3421 0 1000K  
C7310 3421 0 2.5PF   
X734 3520 0 3521 SB 
R7340 3521 0 1000K  
C7340 3521 0 2.5PF   
X737 3620 0 3621 SB 
R7370 3621 0 1000K  
C7370 3621 0 2.5PF   
X740 3720 0 3721 SB 
R7400 3721 0 1000K  
C7400 3721 0 2.5PF   
C7201 2021 0 0.4PF  
C720 2020 0 0.4PF   
C7203 263 0 0.4PF   
C7204 264 0 0.4PF   
L7201 2021 2020 0.1NH       
L7203 263 264 0.1NH 
*   
** OUTPUT IMPEDANC7E
*   
C7MODUL72 264 0 2.5PF       
*********************************************************** 
**************************************************************      
***	8TH ROW 
*********************************************************** 
X81 2050 0 3150 TL  
X82 3150 0 3250 TL  
X83 3250 0 3350 TL  
X84 3350 0 3450 TL  
X85 3450 0 3550 TL  
X86 3550 0 3650 TL  
X87 3650 0 3750 TL  
X88 3750 0 273 TL   
X822 3150 0 3151 SB 
R8220 3151 0 1000K  
C8220 3151 0 2.5PF   
X825 3250 0 3251 SB 
R8250 3251 0 1000K  
C8250 3251 0 2.5PF   
X828 3350 0 3351 SB 
R8280 3351 0 1000K  
C8280 3351 0 2.5PF   
X831 3450 0 3451 SB 
R8310 3451 0 1000K  
C8310 3451 0 2.5PF   
X834 3550 0 3551 SB 
R8340 3551 0 1000K  
C8340 3551 0 2.5PF   
X837 3650 0 3651 SB 
R8370 3651 0 1000K  
C8370 3651 0 2.5PF   
X840 3750 0 3751 SB 
R8400 3751 0 1000K  
C8400 3751 0 2.5PF   
C8201 2051 0 0.4PF  
C820 2050 0 0.4PF   
C8203 273 0 0.4PF   
C8204 274 0 0.4PF   
L8201 2051 2050 0.1NH       
L8203 273 274 0.1NH 
*   
** OUTPUT IMPEDANC8E
*   
C8MODUL82 274 0 2.5PF       
*********************************************************** 
**************************************************************      
*********************************************************** 
*************************************************************** 
*    COLUMN  TL 
*************************************************************** 
XC11 20 0 50 TL     
XC12 1120 0 1150 TL 
XC13 1220 0 1250 TL 
XC14 1320 0 1350 TL 
XC15 1420 0 1450 TL 
XC16 1520 0 1550 TL 
XC17 1620 0 1650 TL 
XC18 1720 0 1750 TL 
XC21 50 0 80 TL     
XC22 1150 0 1180 TL 
XC23 1250 0 1280 TL 
XC24 1350 0 1380 TL 
XC25 1450 0 1480 TL 
XC26 1550 0 1580 TL 
XC27 1650 0 1680 TL 
XC28 1750 0 1780 TL 
XC31 80 0 1020 TL   
XC32 1180 0 2120 TL 
XC33 1280 0 2220 TL 
XC34 1380 0 2320 TL 
XC35 1480 0 2420 TL 
XC36 1580 0 2520 TL 
XC37 1650 0 2620 TL 
XC38 1750 0 2720 TL 
XC41 1020 0 1050 TL 
XC42 2120 0 2150 TL 
XC43 2220 0 2250 TL 
XC44 2320 0 2350 TL 
XC45 2420 0 2450 TL 
XC46 2520 0 2550 TL 
XC47 2620 0 2660 TL 
XC48 2720 0 2750 TL 
XC51 1050 0 1080 TL 
XC52 2150 0 2180 TL 
XC53 2250 0 2280 TL 
XC54 2350 0 2380 TL 
XC55 2450 0 2480 TL 
XC56 2550 0 2580 TL 
XC57 2650 0 2680 TL 
XC58 2750 0 2780 TL 
XC61 1080 0 2020 TL 
XC62 2180 0 3120 TL 
XC63 2280 0 3220 TL 
XC64 2380 0 3320 TL 
XC65 2480 0 3420 TL 
XC66 2580 0 3520 TL 
XC67 2680 0 3620 TL 
XC68 2780 0 3720 TL 
XC71 2020 0 2050 TL 
XC72 3120 0 3150 TL 
XC73 3220 0 3250 TL 
XC74 3320 0 3350 TL 
XC75 3420 0 3450 TL 
XC76 3520 0 3550 TL 
XC77 3620 0 3650 TL 
XC78 3720 0 3750 TL 
.OPTIONS LIMPTS=150000 CPTIME=150000 ITL5=15000 RELTOL=0.001
V2S 201 0 PWL(0.0NS 5 5.2NS 5 5.3NS 0 10.3NS 0 10.4NS 5 15.0NS 5)   
.TRAN 0.03NS 15.0NS UIC     
.PRINT TRAN V(1150) (-5,10) V(51) (-5,10) V(201) (-5,10) V(1281) (-5,10)    
.END
