magic
tech mcnc8
timestamp 641072564
<< polysilicon >>
rect -9 59 -4 63
rect 7 59 40 63
rect -282 31 -276 35
rect -44 31 -39 35
rect -34 20 -29 40
rect 36 40 40 59
rect 55 55 66 59
rect 106 55 109 59
rect 113 55 125 59
rect 136 55 139 59
rect 148 55 156 59
rect 173 55 176 59
rect 186 55 192 59
rect 211 55 214 59
rect -282 16 -276 20
rect -44 16 -39 20
rect -34 16 -10 20
rect 6 16 9 20
rect -34 10 -29 16
rect -34 6 -28 10
rect 23 6 40 10
rect -37 -4 -18 0
rect 12 -4 15 0
rect 36 -17 40 6
rect 51 3 55 48
rect 113 18 117 55
rect 148 30 152 55
rect 186 31 190 55
rect 134 26 152 30
rect 103 14 117 18
rect 51 -1 69 3
rect 77 -1 82 3
rect 148 2 152 26
rect 182 27 190 31
rect 186 2 190 27
rect 114 -2 127 2
rect 138 -2 141 2
rect 148 -2 153 2
rect 179 -2 182 2
rect 186 -2 193 2
rect 212 -2 215 2
rect 114 -17 118 -2
rect 36 -21 118 -17
<< ndiffusion >>
rect -276 -2 -44 16
rect -10 15 6 16
rect -28 10 23 15
rect -28 1 23 6
rect -18 0 12 1
rect -18 -15 -13 -4
rect 69 3 77 4
rect 69 -2 77 -1
<< pdiffusion >>
rect 66 59 106 63
<< metal1 >>
rect 99 74 157 82
rect -40 63 -4 74
rect 7 63 66 74
rect 150 71 157 74
rect 150 70 159 71
rect -40 51 -29 63
rect 109 59 125 70
rect 150 59 156 70
rect 173 59 192 70
rect -286 35 -276 46
rect -11 48 -4 59
rect 7 48 44 59
rect -11 46 6 48
rect -286 31 -279 35
rect -14 31 6 46
rect 66 43 79 44
rect -44 29 -10 31
rect -44 21 -25 29
rect -18 21 -10 29
rect -44 20 -10 21
rect -286 -2 -279 20
rect 36 -2 47 29
rect 69 32 79 43
rect 109 32 117 59
rect 128 33 136 44
rect 69 21 117 32
rect 134 22 136 33
rect 69 15 80 21
rect 92 -2 99 7
rect -286 -13 -276 -2
rect -44 -4 -38 -2
rect 25 -4 69 -2
rect -44 -13 -13 -4
rect -38 -15 -13 -13
rect 12 -13 69 -4
rect 80 -13 99 -2
rect 109 -2 117 21
rect 128 13 136 22
rect 163 31 173 44
rect 163 20 171 31
rect 163 14 173 20
rect 161 13 178 14
rect 201 13 211 44
rect 109 -13 127 -2
rect 152 -13 153 -2
rect 179 -13 193 -2
rect 12 -15 25 -13
rect 92 -17 99 -13
rect 153 -17 159 -13
rect 92 -25 159 -17
rect -368 -103 -103 -39
rect -367 -105 -100 -103
rect -367 -112 -102 -105
rect -367 -114 -100 -112
<< metal2 >>
rect -26 21 -25 28
rect -18 21 -17 28
rect -26 -40 -17 21
rect -103 -105 34 -40
rect -103 -112 -102 -105
rect -94 -112 34 -105
<< polycontact >>
rect -40 40 -29 51
rect -289 20 -278 31
rect 44 48 55 59
rect 36 29 47 40
rect 123 22 134 33
rect 92 7 103 18
rect 171 20 182 31
<< ndcontact >>
rect -276 35 -44 46
rect -276 20 -44 31
rect -10 20 6 31
rect -276 -13 -44 -2
rect -13 -15 12 -4
rect 69 4 80 15
rect 127 2 138 13
rect 153 2 179 13
rect 193 2 212 13
rect 69 -13 80 -2
rect 127 -13 138 -2
rect 153 -13 179 -2
rect 193 -13 212 -2
<< pdcontact >>
rect -4 63 7 74
rect 66 63 106 74
rect 125 59 136 70
rect 156 59 173 70
rect 192 59 211 70
rect -4 48 7 59
rect 66 44 106 55
rect 125 44 136 55
rect 156 44 173 55
rect 192 44 211 55
<< m2contact >>
rect -25 21 -18 29
rect -102 -112 -94 -105
<< ntransistor >>
rect -276 31 -44 35
rect -276 16 -44 20
rect -10 16 6 20
rect -28 6 23 10
rect -18 -4 12 0
rect 69 -1 77 3
rect 127 -2 138 2
rect 153 -2 179 2
rect 193 -2 212 2
<< ptransistor >>
rect -4 59 7 63
rect 66 55 106 59
rect 125 55 136 59
rect 156 55 173 59
rect 192 55 211 59
<< labels >>
rlabel metal1 -10 39 -10 39 1 int
rlabel metal1 -35 68 -35 68 1 Vdd
rlabel metal1 102 26 102 26 1 out
rlabel metal1 167 28 167 28 1 rout
rlabel metal1 36 -10 36 -10 8 GND
rlabel metal1 207 29 207 29 1 load
rlabel polysilicon -36 -2 -36 -2 3 in
<< end >>
