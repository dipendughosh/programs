*Tank anlaysis, ur = 795, sigma = 1.648e5
.OPTIONS ACCT reltol=.0001 abstol=1.0e-15 gmin=1.0e-19
G202B 0 202 102 0 0.1570711544
G202D 0 202 201 0 11.4426022385
G102A 0 102 202 0 0.1111111111
G102C 0 102 103 0 7.7663619448
G201C 0 201 202 0 22.4025140599
G201D 0 201 201 0 85.0762141085
G103D 0 103 102 0 6.5187867813
R102 102 0 0.0514636615
R103 103 0 0.0754159428
R201 201 0 0.0092580181
R202 202 0 0.0506464656
IX302 0 202 AC 0.0000343149 0.0e+00
vtmp 0 5 4
rtmp 5 102 1
.AC LIN 1 60.00 60.00
.WIDTH OUT=80
.PRINT AC VR(102) VR(103) 
.PRINT AC VR(201) VR(202) VR(203) 
.END

