ACTIVE 5TH ORDER LOW-PASS FILTER USING UA741 OPAMP

X0 1 2 ACTIVE
*VIN 1 0 DC 1 AC 1 PULSE( -1 1 )
*VIN 1 0 DC 1 AC 1 PWL( 0 -1 300us -1 330us 1 3.3ms 1 )
VIN 1 0 PWL( 0 -1 300us -1 330us 1 3.3ms 1 )
*wave 1 0 pie { 0,-1 300us,-1 330us,1 3.3ms,1 }

.WIDTH IN=72 OUT=72
.OPT ACCT ITL1=1000 ITL2=1000 ITL5=50000 LIMPTS=1000 reltol=1.0e-6
*.DC VIN -20 20 2
*.AC DEC 25 1 10GHZ
.TRAN 30US 3MS
*.PLOT DC V(2)
*.PLOT AC VM(2)
*.PLOT AC VP(2)
.PRINT TRAN V(1) V(2)

.SUBCKT ACTIVE 100 5
X1 6 0 1 UA741
X2 7 8 2 UA741
X3 9 0 3 UA741
X4 10 11 4 UA741
X5 12 0 5 UA741
C1 6 1 54.63NF
C2 8 0 41.62NF
C3 9 3 106.157NF
C4 11 0 58.79NF
C5 5 12 48.577NF
C13 1 9 26.77NF
C31 6 3 26.77NF
C35 3 12 8.617NF
C53 9 5 8.617NF
R11 6 1 1K
R12 6 100 1K
R13 6 2 1K
R21 7 0 1K
R22 7 2 1K
R23 8 2 1K
R24 8 1 2K
R25 8 3 2K
R31 9 2 1K
R32 9 4 1K
R41 10 0 1K
R42 10 4 1K
R43 11 4 1K
R44 11 3 2K
R45 11 5 2K
R51 12 4 1K
R52 12 5 1K
.ENDS ACTIVE

*.SUBCKT OPAMP 1 2 3
*E0 3 0 2 1 1T
*.ENDS OPAMP

*.SUBCKT SA741 1 2 3
*E1 4 0 2 1 100000
*V1 5 0 13.5V
*V2 0 6 13.5V
*D1 3 5 DIODE
*D2 6 3 DIODE
*R1 1 0 1G
*R2 2 0 1G
*R3 1 2 1MEG
*R4 4 3 100
*C1 3 0 160UF
*.MODEL DIODE D
*.ENDS SA741

.SUBCKT UA741 2 1 24
VCC 27 0 15
VEE 26 0 -15
R1 10 26 1K
R2 9 26 50K
R3 11 26 1K
R4 12 26 3K
R5 15 17 39K
R6 21 20 40K
R7 14 26 50K
R8 18 26 50
R9 24 25 25
R10 23 24 50
R11 13 26 50K
COMP 22 8 30PF
Q1 3 1 4 QML
Q2 3 2 5 QML
Q3 7 6 4 QPL
Q4 8 6 5 QPL
Q5 7 9 10 QML
Q6 8 9 11 QML
Q7 27 7 9 QML
Q8 6 15 12 QML
Q9 15 15 26 QML
Q10 3 3 27 QPL
Q11 6 3 27 QPL
Q12 17 17 27 QPL
Q14 22 17 27 QPL
Q15 22 22 21 QML
Q16 22 21 20 QML
Q17 13 13 26 QML
Q18 27 8 14 QML
Q19 20 14 18 QML
Q20 22 23 24 QML
Q21 13 25 24 QPL
Q22 27 22 23 QML
Q23 26 20 25 QPL
.MODEL QML NPN(BF=80 RB=100 CCS=2PF TF=0.3NS TR=6NS CJE=3PF CJC=2PF
+   VA=50)
.MODEL QPL PNP(BF=10 RB=20 TF=1NS TR=20NS CJE=6PF CJC=4PF VA=50)
.ENDS UA741

.END
