
Rone 4 3 4k
lone 3 0 2m


VIN 4 0 2.5 AC 2.0 0.0
.ac dec 1 1MEG 1MEG
.print ac vp(4) vm(4) vm(4,3) vm(3) vp(3)
.options limpts=10000
.end




