CCSOR CKT - CONSTANT CURRENT SOURCE
*
.MODEL Q1 NPN(BF=49.5 BR=0.5 IS=9.802E-16)

VEE 7 0 -12
VBIAS 3 0 -6.0
Q1 2 3 4 Q1
Q2 2 4 5 Q1
Q3 1 6 5 Q1
Q4 1 8 6 Q1
Q5 10 1 9 Q1
Q6 10 9 8 Q1
R1 2 0 2K
R2 1 0 2K
R3 5 7 2K
R4 8 7 2K
R5 10 0 107


.DC VBIAS -6 6 0.1
.PRINT DC V(1) V(8)
.END
