ECLGATE CKT - ECL STACKED LOGIC GATE

.MODEL D1 D(RS=40 TT=0.1NS CJO=0.9PF)
.MODEL QND NPN(BF=50 RB=70 RC=40 CCS=2PF TF=0.1NS TR=10NS
+ CJE=0.9PF CJC=1.5PF PC=0.85 VA=50)

VEE 15 0 -6.0
VIN 16 0 PULSE(-1.8 -0.8 1NS 1NS 1NS)
VGATE 17 0 PULSE(-0.8 -1.8 5NS 1NS 1NS 5NS)
RS1 16 1 50
Q1 2 1 3 QND
Q2 0 9 3 QND
RC 0 2 100
RS2 17 4 50
Q3 0 4 5 QND
R1 5 6 60
R2 6 15 820
Q4 3 6 7 QND
RE 7 15 280
Q5 0 12 7 QND
R5 0 8 100
Q6 0 8 9 QND
R3 9 15 2K
D1 8 10 D1
R6 10 11 60
Q7 0 11 12 QND
R4 12 15 2K
D2 11 13 D1
R7 13 15 720
Q8 0 2 14 QND
RL 14 15 560


.TRAN 0.1NS 20NS
.PRINT TRAN V(16) V(17) V(6) V(14)
.END

