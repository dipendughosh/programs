
G102A 0 102 202 0 1.0
G102C 0 102 103 0 2.0

R102 102 0 0.05
R103 103 0 0.07
R105 103 202 70

R202 202 0 0.05

IX302 0 202 0.0 AC 0.00003 0.0e+00

.OPTIONS ACCT reltol=.0001 abstol=1.0e-15 gmin=1.0e-19
.AC LIN 1 60.00 60.00
.WIDTH OUT=80
.PRINT AC VR(102) VR(202) 
.END

