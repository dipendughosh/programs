256 DRAM CONTROL CHAIN CIRCUIT 
*****************************************************
*     N-CHANNEL LOW ENHANCEMENT TRANSISTOR MODEL  *
*****************************************************
.MODEL ML NMOS LEVEL=3
+ RSH=0 TOX=300e-10 LD=0.21e-6 XJ=0.28e-6 VMAX=15e4 ETA=0.18
+ KAPPA=0.5 NSUB=2.8e14 UO=730 THETA=0.095 VTO=0.5 CGSO=2.8e-10
+ CGDO=2.8e-10 CJ=5.7e-5 CJSW=2.48e-10 PB=0.7 MJ=0.5 MJSW=0.3
+ NFS=1e10

*****************************************************
*     N-CHANNEL HIGH ENHANCEMENT TRANSISTOR MODEL *
*****************************************************
.MODEL MH NMOS LEVEL=3
+ RSH=0 TOX=300e-10 LD=0.21e-6 XJ=0.28e-6 VMAX=15e4 ETA=0.18
+ KAPPA=0.5 NSUB=3.5e14 UO=700 THETA=0.095 VTO=0.8 CGSO=2.8e-10
+ CGDO=2.8e-10 CJ=5.7e-5 CJSW=2.48e-10 PB=0.7 MJ=0.5 MJSW=0.3
+ NFS=1e10

*****************************************************
*     N-CHANNEL DEPLETION TRANSISTOR MODEL        *
*****************************************************
.MODEL MD NMOS LEVEL=3
+ RSH=0 TOX=300e-10 LD=0.21e-6 XJ=0.28e-6 VMAX=15e4 ETA=0.18
+ KAPPA=0.5 NSUB=3.5e14 UO=700 THETA=0.035 VTO=-3.0 CGSO=2.8e-10
+ CGDO=2.8e-10 CJ=5.7e-5 CJSW=2.48e-10 PB=0.7 MJ=0.5 MJSW=0.3
+ NFS=1e10


*****************************
* PAGE 1
*****************************


* SIMULATION CIRCUIT ITEMS
CCRE     11  0 2p
CCRE1     12  0 2p
CNCRE     778 0 1p
CCER     51  0 3p
CCE1R     52  0 3p
CPCRTR     54  0 2.8p
CCERN     251 0 0.63p
CCE1RN     252 0 0.63p
CPCRTRN     254 0 1.03p
CCCDE     59  0 2p
CPCDB     57  0 2p
CPCDBP     58  0 1p
CCCEL     56  0 2p
CPRDB     14  0 1p
CPRDBP     15  0 1p

* CIRCUIT BLOCK

M118     1     1     107 9999 ML W=5U   L=2U
M119     1     104     107 9999 MH W=5U   L=2U
M121     107     104     108 9999 ML W=15U  L=2U
M123     108     104     109 9999 MH W=15U  L=2U
M125     109     13     0   9999 MH W=17U  L=2U
M130     1      13     108 9999 MH W=2U   L=3U
M122     1     107     103 9999 MH W=140U L=2U
M111     1      1     103 9999 ML W=44U  L=2U
M106     103     103     104 9999 MD W=3.5U L=15U
M108     104     10     110 9999 ML W=200U L=2U
M128     110     10     0   9999 MH W=250U L=2U
M126     1     104     110 9999 MH W=7U   L=2U
M109     1     104     11  9999 MH W=215U L=2U
M110     11     10     0   9999 MH W=100U L=2.5U
M112     11     103     11  9999 MD W=200U L=60U
M113     1     11     12  9999 ML W=100U L=2.25U
M114     12     10     0   9999 MH W=75U  L=2.5U
M124     15     107     15  9999 MH W=20U  L=20U

*****************************
* PAGE 2
*****************************

M162     1     155     155 9999 MH W=5U    L=2U
M163     155     154     154 9999 MH W=5U    L=2U
M161     1     1     154 9999 ML W=15U   L=2U
M166     154     10     156 9999 MH W=60U   L=3U
M167     156     10     157 9999 MH W=40U   L=2U
M168     157     11     0   9999 MH W=40U   L=2U
M165     1     154     156 9999 MH W=3U    L=2U
M164     11     154     11  9999 MH W=15U   L=20U
M158     1     11     152 9999 ML W=15U   L=2.25U
M159     152     10     0   9999 MH W=50U   L=2U
M160     1     154     151 9999 ML W=70U   L=2U
M169     151     151     1511 9999 MD W=3U   L=15U
M155     1511     152     153 9999 MH W=60U   L=2U
M156     153     152     0   9999 MH W=60U   L=2U
M157     1     1511     153 9999 MH W=3U    L=2U
M154     150     151     150 9999 MD W=400U  L=3U
M152     1     1511     150 9999 ML W=50U   L=2.25U
M153     150     12     0   9999 MH W=20U   L=2U
M150     1     1511     13  9999 ML W=400U  L=2.25U
M151     13     12     0   9999 MH W=500U  L=2U

******************************
* NEW CRE DELAY BLOCK
******************************
M711     1     1     703 9999 ML W=20U  L=2U
M703     703     703     704 9999 MD W=3.5U  L=10U
M708     704     777     710 9999 ML W=5U  L=2U
M728     710     777     0   9999 MH W=5U  L=2U
M726     1     704     710 9999 MH W=3U  L=2U
M709     1     704     778 9999 MH W=100U  L=2U
M710     778     777     0   9999 MH W=50U  L=2U
M712     778     703     778 9999 MD W=20U  L=10U
M713     1     13     777 9999 ML W=20U  L=2U
M714     777     11     0   9999 MD W=40U  L=2U

******************************
* CIRCUIT BLOCK (PRDB & PRDBP BLOCK)
******************************

M5141     1     504     504 9999 ML W=20U  L=2U
M514      1     1     504 9999 ML W=10U  L=2U
M510      13     504     13  9999 MH W=10U  L=5U
M513      13     504     5011 9999 ML W=100U  L=2U
M515      504     1     5041 9999 ML W=15U  L=2U
M522      5041     509     506 9999 ML W=15U  L=2U
M523      506     11     0   9999 MH W=10U  L=2U

M524      0     506     0   9999 MD W=10U  L=10U
M516      5011     1     507 9999 MH W=15U  L=2U
M517      507     11     0   9999 MH W=15U  L=2U
M505      5011     5011     501 9999 MD W=3U  L=15U
M504      509     5011     509 9999 MD W=100U  L=10U
M511      1     13     503 9999 MH W=6U  L=3U
M512      503     11     0   9999 ML W=10U  L=2.25U
M500      1     11     502 9999 ML W=20U  L=2.25U
M593      502     503     0   9999 MH W=20U  L=3U
M506      501     502     505 9999 MH W=80U  L=2U
M508      505     502     0   9999 MH W=100U  L=2U
M507      1     501     505 9999 MH W=3U  L=2U
M527      508     501     509 9999 ML W=50U  L=2.25U
M528      508     501     14  9999 MH W=200U  L=2.25U
M509      509     502     505 9999 MH W=100U  L=2U
M533      1     1     14  9999 ML W=2U  L=3U
M530      1     14     531 9999 MH W=4U  L=2U
M531      14     12     531 9999 MH W=400U  L=2U
M532     531     12     0   9999 MH W=400U L=2U

*****************************
* PAGE 3
*****************************
m590 1 11 512 9999 ML w=5u l=2.25u
m501 17 512 511 9999 ML w=30u l=2u
m502 512 1 5121 9999 MH w=5u l=2u
m503 5121 13 0 9999 MH w=5u l=2u
m538 511 15 0 9999 MH w=10u l=2u
m518 511 510 511 9999 MH w=50u l=10u
m519 1 14 510 9999 MH w=10u l=2u
m520 1 1 510 9999 ML w=10u l=2u
m521 510 511 522 9999 MH w=30u l=2u
m525 1 510 508 9999 ML w=200u l=2u
m526 1 1 508 9999 ML W=50u l=2u
m529 15 508 15 9999 ML w=700u l=20u

*PRDBP BLOCK
m544 1 11 524 9999 ML w=5u l=2.25u
m5441 1 524 524 9999 ML w=15u l=2u
m545 13 524 5211 9999 ML w=60u l=2u
m548 524 1 526 9999 MH w=15u l=2u
m549 526 520 0 9999 ML w=15u l=2u
m546 5211 1 527 9999 MH w=15u l=2u
m547 527 11 0 9999 MH w=15u l=2u
m535 5211 5211 521 9999 MD w=3u l=15u
m534 520 5211 520 9999 MD w=100u l=7u
m541 1 14 523 9999 MH w=5u l=3u
m542 523 11 0 9999 MH w=5u l=2u
m539 1 11 522 9999 ML w=20u l=2.25u
m540 522 523 0 9999 MH w=30u l=3u
m550 521 522 525 9999 MH w=70u l=2u
m551 525 522 0 9999 MH w=70u l=2u
m552 1 521 525 9999 MH w=3u l=2u
m553 1 521 520 9999 ML w=20u l=2.25u
m555 1 521 15 9999 ML w=90u l=2u
m554 520 522 0 9999 MH w=20u l=2u
m556 15 528 0 9999 MH w=200u l=2u
m557 1  11 528 9999 ML w=20u l=2.25u
m558 528 13 0 9999 MH w=10u l=2u
rPRDBP 1 15 50k

m3059 1 14 3054 9999 MH w=5u l=2u
m3060 1 3054 3054 9999 ML w=30u l=2u
m3058 1 30511 3054 9999 MH w=10u l=2u
m3061 54 3054 54 9999 MH w=50u l=2u
m3057 17 3054  30511 9999 ML w=100u l=2u
m30621 1 3054 30541 9999 MH w=2u l=3u
m30641 3054 1 30542 9999 MH w=20u l=2u
m3064 30542 0 0  9999 MH w=20u l=2u
m3062 3054 3050 30541 9999 ML w=20u l=2u
m3063  30541 3050 3055 9999 ML w=20u l=2u
m3066 0 3055 0 9999 MD w=75u l=2u
m3065 3055 54 0 9999 ML w=10u l=2u
m3056 3050 30511 3050 9999 MD w=200u l=5u
m3068 30511 1 3056 9999 MH w=15u l=2u
m3069 3056 0 0  9999 ML w=15u l=2u
m3070 3056 13 0 9999 ML w=15u l=2u
m3067 30511 30511 3051 9999 MD w=3u l=15u
m3079 1 17 3053 9999 MH w=5u l=2.5u
m3080 3053 13 0 9999 ML w=5u l=2u
m3077 1 13 3052 9999 ML w=30u l=2u
m3076 1 14 3052 9999 MH w=10u l=2u
m3078 3052 3053 0 9999 MH w=20u l=2.5u
m3075 1 3051 3057 9999 MH w=6u l=2u
m3074 3057 50 0 9999 MH w=100u l=2u
m3073 3057 3052 0 9999 MH w=50u l=2u
m3072 3051 50 3057 9999 MH w=100u l=2u
m3071 3051 3052 3057 9999 MH w=50u l=2u
m3052 1 3051 3050 9999 ML w=30U l=2.25u

*****************************
* PAGE 4
*****************************
m3050 1 3051 51 9999 ML w=300u l=2.25u
m3055 3050 50 0 9999 MH w=30u l=2.5u
m3053 3050 3052 0 9999 MH w=30u l=2u
m3051 51 3052 0 9999 MH w=50u l=2u
m3054 51 50 0 9999 MH w=250u l=2.5u
m3081 51 0 0 9999 MH w=10u l=2u
m3082 51 13 0 9999 ML w=30u l=2u

*CCE1R BLOCK
m3085 1 51 52 9999 MH w=200u l=2u
m3086 52 50 0 9999 MH w=150u l=2.5u
m3088 52 13 0 9999 MH w=30u l=2u
m3095 52 3052 0 9999 MH w=50u l=2u

*CIRCUIT BLOCK (PCRTR & PCRTR1 BLOCK) 
m3214 1 3207 3207 9999 MH w=5u l=2u
m3215 3207 3204 3204 9999 MH w=5u l=2u
m3213 1 1 3204 9999 ML w=15u l=2u
m3205 1 3204 32011 9999 ML w=70u l=2u
m3216 51 3204 51 9999 MH w=100u l=3u
m3212 32011 32011 3201 9999 MD w=3u l=15u
m3204 3203 32011 3203 9999 MD w=70u l=20u
m3219 3204 50 3208 9999 MH w=40u l=2u
m3220 3208 50 3200 9999 MH w=40u l=2u
m3222 3200 51 0 9999 MH w=40u l=2u
m3221 1 3204 3208 9999 MH w=3u l=2u
m3217 3204 1 32041 9999 MH w=10u l=2u
m3218 32041 13 3200 9999 MH w=10u l=2u
m3209 1 51 3202 9999 ML w=6u l=2.25u
m3210 3202 50 0 9999 MH w=50u l=2.5u
m3211 3202 13 0 9999 MH w=30u l=2u
m3206 3201 3202 3233 9999 MH w=60u l=2u
m3207 3233 3202 0 9999 MH w=60u l=2u
m3239 1 3201 3233 9999 MH w=3u l=2u
m3202 1 3201 3203 9999 ML w=50u l=2.25u
m3203 3203 52 0 9999 MH w=50u l=2u
m3223 3201 3203 3223 9999 MH w=20u l=2u
m3224 3223 51 0 9999 MH w=20u l=2u
m3200 1 3201 54 9999 ML w=400u l=2.25u
m3201 54 52 0 9999 MH w=500u l=2u
RPCRTR 1 54 40k

* PCRTR1 BLOCK
m3290 1 54 55 9999 MH w=30u l=2u
m3291 55 51 0 9999 MH w=160u l=2u

* CIRCUIT BLOCK (NEW CCER & CCE1R BLOCK)
m2059 1 14 2054 9999 MH w=5u l=2u
m2060 1 2054 2054 9999 ML w=15u l=2u
m2058 1 20511 2054 9999 MH w=10u l=2u
m2061 254 2054 254 9999 MH w=25u l=2u
m2057 17 2054 20511 9999 ML w=50u l=2u
m20621 1 2054 20541 9999 MH w=2u l=3u
m20641 2054 1 20542 9999 MH w=10u l=2u
m2064 20542 0 0 9999 MH w=10u l=2u
m2062 2054 2050 20541 9999 ML w=10u l=2u
m2063 20541 2050 2055 9999 ML w=10u l=2u
m2066 0 2055 0 9999 MD w=40u l=2u
m2065 2055 254 0 9999 MH w=5u l=2u
m2056 2050 20511 2050 9999 MD w=60u l=5u
m2068 20511 1 2056 9999 MH w=8u l=2u
m2069 2056 0 0 9999 MH w=8u l=2u
m2070 2056 13 0 9999 MH w=8u l=2u
m2067 20511 20511 2051 9999 MD w=3u l=15u
m2079 1 17 2053 9999 MH w=5u l=2.5u
m2080 2053 13 0 9999 MH w=5u l=2u

*****************************
* PAGE 5
*****************************

m2077     1    13  2052  9999 ML W= 13u L= 2u
m2076     1    14  2052  9999 MH W=  5u L= 2u
m2078  2052  2053     0  9999 MH W= 10u L= 2.5u
m2075     1  2051  2057  9999 MH W=  3u L= 2u
m2074  2057    50     0  9999 MH W= 50u L= 2u
m2073  2057  2052     0  9999 MH W= 25u L= 2u
m2072  2051    50  2057  9999 MH W= 50u L= 2u
m2071  2051  2052  2057  9999 MH W= 25u L= 2u
m2052     1  2051  2050  9999 ML W= 15u L= 2.25u
m2050     1  2051   251  9999 ML W=100u L= 2.25u
m2055  2050    50     0  9999 MH W= 10u L= 2.5u
m2053  2050  2052     0  9999 MH W= 15u L= 2u
m2051   251  2052     0  9999 MH W= 25u L= 2u
m2054   251    50     0  9999 MH W= 80u L= 2.5u
m2081   251     0     0  9999 MH W=  5u L= 2u
m2082   251    13     0  9999 MH W= 15u L= 2u

*CCE1R BLOCK
m2085     1   251   252  9999 MH W= 50u L= 2u
m2086   252    50     0  9999 MH W= 40u L= 2.5u
m2088   252    13     0  9999 MH W= 10u L= 2u
m2095   252  2052     0  9999 MH W= 15u L= 2u

* CIRCUIT BLOCK (NEW PCRTR BLOCK)
m2214     1  2207  2207  9999 MH W=  5u L= 2u
m2215  2207  2204  2204  9999 MH W=  5u L= 2u
m2213     1     1  2204  9999 ML W= 15u L= 2u
m2205     1  2204 22011  9999 ML W= 35u L= 2u
m2216   251  2204   251  9999 MH W= 50u L= 3u
m2212 22011 22011  2201  9999 MD W=  3u L=15u
m2204  2203 22011  2203  9999 MD W= 70u L=10u
m2219  2204    50  2208  9999 MH W= 40u L= 2u
m2220  2208    50  2200  9999 MH W= 40u L= 2u
m2222  2200   251     0  9999 MH W= 40u L= 2u
m2221     1  2204  2208  9999 MH W=  3u L= 2u
m2217  2204     1 22041  9999 MH W= 10u L= 2u
m2218 22041    13  2200  9999 MH W= 10u L= 2u
m2209     1   251  2202  9999 ML W=  4u L= 2.25u
m2210  2202    50     0  9999 MH W= 25u L= 2.5u
m2211  2202    13     0  9999 MH W= 15u L= 2u
m2206  2201  2202  2233  9999 MH W= 30u L= 2u
m2207  2233  2202     0  9999 MH W= 30u L= 2u
m2239     1  2201  2233  9999 MH W=  3u L= 2u
m2202     1  2201  2203  9999 ML W= 25u L= 2.25u
m2203  2203   252     0  9999 MH W= 25u L= 2u
m2223  2201  2203  2223  9999 MH W= 10u L= 2u
m2224  2223   251     0  9999 MH W= 10u L= 2u
m2200     1  2201   254  9999 ML W=200u L= 2.25u
m2201   254   252     0  9999 MH W=300u L= 2u
RPCRTRN   1   254   40K

* CIRCUIT BLOCK (CCDE BLOCK)
m1117     1    54  1104  9999 ML W= 20u L= 2u
m1116     1  1104  1104  9999 ML W= 30u L= 2u
m1106    51  1104  1105  9999 ML W=150u L= 2u
m1105  1105  1104 11011  9999 ML W=150u L= 2u
m1118     1 11011  1105  9999 MH W=  3u L= 2u
m1119  1104     1 11041  9999 MH W= 30u L= 2u
m1120 11041  1100     0  9999 ML W= 30u L= 2.25u
m1104  1100 11011  1100  9999 MD W= 60u L=20u
m1115 11011 11011  1101  9999 MD W=  3u L=13u
m1113     1    51  1103  9999 MH W= 15u L= 3u
m1114  1103    54     0  9999 MH W= 15u L= 2u
m1110     1    51  1102  9999 ML W= 30u L= 2u
m1111     1    14  1102  9999 MH W= 10u L= 2u
m1112  1102  1103     0  9999 MH W= 50u L= 2.3u

*****************************
* PAGE 6
*****************************

m1107 1101 1102 1106 9999 ML w=60u l=20u
m1109 1 1101 1106 9999 MH w=3u l=2u
m1108 1106 1102 0 9999 MH w=60u l=2u
m1102 1 1101 1100 9999 ML w=50u l=2.25u
m1103 1100 1102 0 9999 MH w=50u l=2u
m1100 1 1101 59 9999 ML w=400u l=2.25u
m1101 59 1102 0 9999 MH w=250u l=2u

* CIRCUIT BLOCK (PCDB BLOCK)
m1394 1 1307 1307 9999 MH w=10u l=2u
m1395 1 1 1307 9999 ML w=10u l=2u
m1322 1 59 1304 9999 ML w=10u l=2.25u
m1323 1 1304 1304 9999 ML w=15u l=2.25u
m1320 54 1304 1303 9999 ML w=170u l=2u
m1321 1 13011 1303 9999 MH w=3u l=2u
m1324 1304 1 13041 9999 MH w=20u l=2u
m1325 13041 1300 0 9999 ML w=20u l=2u
m1319 1303 1307 13011 9999 ML w=170u l=2u
m1396 1307 1 13071 9999 MH w=20u l=2u
m1397 13071 1300 1305 9999 ML w=20u l=2u
m1326 0 1305 0 9999 MD w=10u l=30u
m1327 1305 59 0 9999 MH w=10u l=2u
m1310 1300 13011 1300 9999 MD w=100u l=20u
m1311 13011 13011 1301 9999 MD w=3u l=10u
m1335 1 51 1313 9999 ML w=5u l=2.25u
m1336 61 1313 1312 9999 ML w=30u l=2u
m1337 1313 1 13131 9999 MH w=5u l=2u
m1338 13131 54 0 9999 MH w=5u l=2u
m1339 1312 58 0 9999 MD w=10u l=2u
m1399 1 59 1302 9999 MH w=5u l=2u
m1334 1312 1311 1312 9999 MH w=50u l=10u
m1333 1311 1312 1322 9999 MH w=30u l=2u
m1331 1 57 1311 9999 MH w=10u l=2u
m1332 1 1 1311 9999 ML w=10u l=2u
m1330 1 1311 1310 9999 ML w=250u l=2u
m1329 1 1 1310 9999 ML w=50u l=2u
m1328 58 1310 58 9999 ML w=800u l=20u
m1317 1 54 1309 9999 MH w=6u l=2u
m1318 1309 59 0 9999 MH w=5u l=2u
m13181 1309 51 0 9999 MH w=5u l=2u
m1315 1 51 1302 9999 ML w=30u l=2.25u
m1316 1302 1309 0 9999 MH w=30u l=2u
m1312 1301 1302 1306 9999 MH w=100u l=2u
m1314 1 1301 1306 9999 MH w=3u l=2u
m1313 1306 1302 0 9999 MH w=150u l=2u
m1306 1310 1301 1300 9999 ML w=60u l=2.25u
m1300 1310 1301 57 9999 ML w=250u l=2.25u
m1340 1 1 57 9999 ML w=3u l=30u
m1305 1 57 1308 9999 MH w=4u l=2u
m1304 1308 52 0 9999 MH w=400u l=2u
m1303 57 52 1308 9999 MH w=400u l=2u
m1307 1300 1302 1306 9999 MH w=100u l=2u
m1301 57 1302 1306 9999 MH w=50u l=2u

* PCDB BLOCK
m1383 1 59 1324 9999 ML w=10u l=2.25u
m1384 1 1324 1324 9999 ML w=15u l=2.25u
m1381 54 1324 1326 9999 ML w=100u l=2u
m1385 1324 1 13241 9999 MH w=15u l=2u
m1386 13241 1320 0 9999 ML w=15u l=2u
m1382 1 13211 1326 9999 MH w=3u l=2u
m1380 1326 1324 13211 9999 ML w=100u l=2u
m1374 1320 13211 1320 9999 MD w=70u l=10u
m1375 13211 13211 1321 9999 MD w=3u l=15u
m1387 54 57 1323 9999 MH w=5u l=2u
m1388 1323 59 0 9999 MH w=5u l=2u



*****************************
* PAGE 7
*****************************
M1389     1     51     1322   9999 ML w=20u l=2.25u
M1390     1322     1323     0      9999 MH w=20u l=2u
M1391     1     59     1322   9999 MH w=5u l=2u
M1377     1321     1322     1325   9999 MH w=3u l=2u
M1378     1325     1322     0      9999 MH w=70u l=2u
M1379     1     1321     1325   9999 MH w=3u l=2u
M1372     1     1321     1320   9999 ML w=25u l=2.25u
M1371     1321     1320     13212  9999 MH w=20u l=2u
M1392     13212     51     0      9999 MH w=20u l=2u
M1373     1320     1322     0      9999 MH w=25u l=2u
M1370     1     1321     58     9999 ML w=100u l=2.25u
M1393     1     1     58     9999 ML w=3u l=30u
M1398     58     1302     0      9999 MH w=25u l=2u
M1376     58     52     0      9999 MH w=200u l=2u

* CIRCUIT BLOCK (CCEL BLOCK)
M1064     1     14     1054     9999 MH w=5u l=2u
M1065     1     1054     1054     9999 ML w=30u l=2u
M1066     1     10511     1054     9999 MH w=10u l=2u
M1067     57     1054     57     9999 MH w=10u l=10u
M10661     1     1054     10541     9999 MH w=2u l=3u
M1055     17     1054     10511     9999 ML w=100u l=2u
M1068     1054     1050     10541     9999 ML w=20u l=2u
M1069     10541     1050     1055     9999 ML w=20u l=2u
M1072     0     1055     0     9999 MD w=75u l=2u
M1071     1055     57     0     9999 MH w=20u l=2u
M1054     1050     10511     1050     9999 MD w=100u l=10u
M1056     10511     10511     1051     9999 MD w=3u l=15u
M1060     1     57     1056     9999 MH w=10u l=2u
M1061     55     1056     55     9999 MH w=20u l=3u
M1062     1056     59     0     9999 MH w=5u l=3u
M1063     1     13     55     9999 ML w=30u l=2u
M1057     1051     55     1053     9999 MH w=70u l=2u
M1059     1     1051     1053     9999 MH w=3u l=2u
M1058     1053     55     0     9999 MH w=70u l=2u
M1052     1     1051     1050     9999 ML w=25u l=2.25u
M1073     1051     1050     11     9999 MH w=20u l=2u
M1050     1     1051     56     9999 ML w=250u l=2.25u
M1053     1050     55     0     9999 MH w=25u l=2u
M1051     56     55     0     9999 MH w=200u l=2u

.options nopage nomod limpts=100000 itl1=500 itl5=100000 reltol=0.01
.width in=80 out=132
.print tran v(51) v(52) v(50) v(54) v(55) v(56) v(251) v(252) v(254)
+  v(58) v(59) v(61)
.print tran v(10) v(11) v(12) v(13) v(17) v(778) v(14) v(15)

.ic v(10)=3v v(11)=0v v(12)=0v v(13)=5v v(17)=0v v(54)=0v v(14)=5v
+   v(50)=3v v(51)=0v v(52)=0v v(59)=5v v(58)=5v v(57)=8v v(61)=0v
+   v(56)=0v v(15)=5v v(251)=0v v(252)0v v(254)=5v

* VOLTAGE SOURCES
VCC 1 0 DC 5V
VBB 0 9999 DC 2.5V
VRE 10 0     PWL(0 3.0v 5n 3.0V 8n 0.0v 110n 0.0v 113n 3.0v 120n 3.0v)
VCR 17 0     PWL(0 0.0v 30n 0.0v 35n 5.0v 120n 5v)
VCE 50 0     PWL(0 3.0v 50n 3.0v 53n 0.0v 105n 0.0v 108n 3.0v 120n 3.0v)
VCCAV 61 0     PWL(0 0.0v 75n 0.0v 80n 5.0v 120n 5v)

.tran 0.1ns 120ns
.end
