
Rone 4 3 10k
Cone 3 0 2p


VIN 4 0 2.5 AC 2.0 0.0
.ac dec 10 1MEG 10000MEG
.print ac ir(VIN) ii(VIN)
.options limpts=10000
.end



