CFFLOP CKT - SATURATING COMPLEMEMTARY FLIP-FLOP

.MODEL QN1 NPN(BF=10 BR=1 IS=9.1E-15)
.MODEL QP1 PNP(BF=10 BR=1 IS=9.1E-15)

VCC1 1 0 5.0
VCC2 8 0 10.0
VEE1 10 0 -5.0
VEE2 9 0 -10.0
Q1 3 2 1 QP1
Q2 6 7 1 QP1
Q3 6 5 10 QN1
Q4 3 4 10 QN1
R1 8 2 57.2K
R2 8 7 57.2K
R3 2 6 14.3K
R4 7 3 14.3K
R5 6 4 14.3K
R6 3 5 14.3K
R7 4 9 57.2K
R8 5 9 57.2K
R9 3 0 1K


CIN 3 99 1U
*VIN 99 0 PULSE(0 1 10NS 20NS 20NS 500NS 1000NS) 
VIN 99 0 SIN(0 1 2MEG 20NS 0 ) 
.TRAN 1NS 1000NS 
.PRINT TRAN V(99) V(3) V(6)
.OPTIONS NUMDGT=6 LIMPTS=10000
.END
