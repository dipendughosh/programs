*** simple inverter for CAzM GaAs verification ***

* typical typical models

.model mfet15 njf 
+ vto=-0.460 beta=2.72e-04 rsh=765 gamds=-0.006 is=3.88e-2 n=1.210 ldel=-0.385u
+ vgexp=2.55 alpha=3.94 ucrit=0.051 lambda=0.127 satexp=3.68
+ ng=0.595 nd=0.100 k1=0.204 eg=876e-03 gap1=1e-06 gap2=10 d=13.1 
+ gcap=1.495e-03 crat=.1109
+ level=3 capop=1 sat=3
+ acm=1 hdif=2.615u rshl=0 rs=0 rd=0 xti=2 tlev=2 
+ trs=2.24e-03 trd=2.24e-03 bex=481e-03 tcv=290e-06

.model mfet04 njf 
+ vto=0.227 beta=3.02e-04 rsh=2171 gamds=-0.041 is=1.02e-2 n=1.227 ldel=-0.385u
+ vgexp=2.35 alpha=6.53 ucrit=1e-4 lambda=0.072 satexp=3.29
+ ng=0.961 nd=0.100 k1=0.224 eg=917e-03 gap1=1e-06 gap2=10 d=13.1
+ gcap=1.062e-03 crat=.1109
+ level=3 capop=1 sat=3
+ acm=1 hdif=0.815u rshl=0 rs=0 rd=0 xti=2 tlev=2 
+ trs=-1.17e-03 trd=-1.17e-03 bex=-2 tcv=1.64e-03

jm1 dm1 gm1 sm1 bm1 mfet04 w=50u l=5u
jm2 dm2 gm2 sm2 bm2 mfet15 w=5u  l=5u

vdm1 dm1 0 2.0
vgm1 gm1 0 2.0
vsm1 sm1 0 2.0
vbm1 bm1 0 2.0

vdm2 dm2 0 2.0
vgm2 gm2 0 2.0
vsm2 sm2 0 2.0
vbm2 bm2 0 2.0

.dc vdm1 0.0 2.0 0.04 vgm1 0.0 0.5 0.1
.print dc lx9(jm1) lx11(jm1) lx13(jm1) lx14(jm1)
.options dccap ingold=2
.end
