
*.model nenh nmos
*+    Level=2            Ld=0.042u       Tox=197.000e-10
*+    Nsub=1.066e+16     Vto=0.381       Kp=1.1601e-04
*+    Gamma=.639243      Phi=.31         Uo=1957.00
*+    Uexp=4.612355e-2   Ucrit=174667    Delta=0.0
*+    Vmax=177269        Xj=.9u          Lambda=0.0
*+    Nfs=4.55168e+12    Neff=4.68830    Nss=3.000000E+10
*+    Tpg=1.00000        Rsh=60          Cgso=2.89e-10
*+    Cgdo=2.89e-10      Cj=3.27e-04     Mj=1.067
*+    Cjsw=1.74e-10      Mjsw=.195

*.model penh pmos
*+    Level=2            Ld=.197u        Tox=209.000e-10  
*+    Nsub=6.575441e+16  Vto=-0.472      Kp=3.816E-05
*+    Gamma=0.618101     Phi=.541111     Uo=488.0
*+    Uexp=8.886957e-02  Ucrit=637449    Delta=0.0
*+    Vmax=63253.3       Xj=0.112799u    Lambda=0.    
*+    Nfs=1.668437e+11   Neff=0.64354    Nss=3.000000E+10
*+    Tpg=-1.00000       Rsh=150         Cgso=3.35e-10
*+    Cgdo=3.35e-10      Cj=4.75e-04     Mj=.341
*+    Cjsw=2.23e-10      Mjsw=.307

*
*
*
.SUBCKT INVERT1 1 2 3 4
.MODEL MOD1 PMOS LEVEL=1  VTO=-0.47 KP=3.816E-05 PHI=0.5411 GAMMA=0.62 
.MODEL MOD2 NMOS LEVEL=1  VTO=0.38  KP=1.1601E-04 PHI=0.31 GAMMA=0.64 
mtwo 2 1 3 3 MOD1 l=1.0u w=1200.0u ad=1200.0p pd=1202.0u as=1200.0p ps=1202.0u
mone 2 1 4 4 MOD2 l=1.0u w=800.0u ad=800.0p pd=802.0u as=800.0p ps=802.0u
.ENDS INVERT1
.SUBCKT INVERT2 1 2 3 4
.MODEL MOD1 PMOS LEVEL=1  VTO=-0.47 KP=3.816E-05 PHI=0.5411 GAMMA=0.62 
.MODEL MOD2 NMOS LEVEL=1  VTO=0.38  KP=1.1601E-04 PHI=0.31 GAMMA=0.64 
mtwo 2 1 3 3 MOD1 l=1.0u w=40.0u ad=40.0p pd=42.0u as=40.0p ps=42.0u
mone 2 1 4 4 MOD2 l=1.0u w=20.0u ad=20.0p pd=22.0u as=20.0p ps=22.0u
.ENDS INVERT2
R1 10 103 0.01
R2 20 203 0.01
R3 30 303 0.01
X11 100 101 88 0 INVERT1
X12 104 105 88 0 INVERT2
X13 200 201 888 0 INVERT1
X14 2044 205 88 0 INVERT2
X15 300 301 88 0 INVERT1
X16 304 305 88 0 INVERT2
C101 101 0 0.4P
C10 10 0 0.4P
C103 103 0 0.4P
C104 104 0 0.4P
C105 105 0 0.1P
L101 101 10 0.1N
L103 103 104 0.1N
C201 2011 0 0.4P
C20 20 0 0.4P
C203 203 0 0.4P
C204 204 0 0.4P
C205 205 0 0.1P
L201 2011 20 0.1N
L203 203 204 0.1N
C301 301 0 0.4P
C30 30 0 0.4P
C303 303 0 0.4P
C304 304 0 0.4P
C305 305 0 0.1P
L301 301 30 0.1N
L303 303 304 0.1N
R103 103 0 100
R203 203 0 100
R303 303 0 100
.OPTIONS LIMPTS=100000 CPTIME=100000 ITL5=100000 RELTOL=0.01
.IC V(100)=3 V(101)=0 V(200)=0 V(201)=3 V(300)=3 V(301)=0
V1S 100 0 DC 3
V3S 300 0 DC 3
VDD 88  0 DC 3
VI88 88 888
VI201 201 2011
VI204 204 2044
V2S 200 0 PWL(0.0NS 0 1NS 3 5NS 3 6NS 0 10NS 0 11NS 3 15NS 3
+16NS 0 20NS 0 21NS 3 25NS 3 26NS 0
+30NS 0 31NS 3 35NS 3 36NS 0 40NS 0)
.TRAN 0.010NS 40NS UIC
*.PRINT TRAN   V(103) V(203) V(303)
.PRINT TRAN  V(88) I(VI88) V(201) I(VI201) V(204) I(VI204)
.END
