* Project TRY1
* WorkVIEW Wirelist Created with Version 4.1

CINT     N56 N57 200P
C1       N20 N56 2.0U
C2       N57 N22 2.0U
L1       N57 N56 200U
R1       N27 0   1K
CEXT     N56 N57 2U
XT1      N56 N57 N27 0   TRANSF
R3       N6  N56 1.0
R2       N8  N57 1.0

* DICTIONARY 8
* $1N27 = N27
* $1N8 = N8
* $1N6 = N6
* $1N22 = N22
* $1N20 = N20
* $1N57 = N57
* $1N56 = N56
* GND = 0
* PROBES 1
* V(N27)


* MODEL FILE FOR "TRANSF" TRANSFORMER SYMBOL
*
* To change the parameters of the transformer, copy this 
* model file to another file and perform the following steps:
*
*		1)	Change the name of the subckt from "TRANSF" to
*			the same name as your file.
*		2)	Change the value of the primary inductance.
*		3)	Change the value of the secondary inductance.
*		4)	Change the coefficient of coupling.
*		5)	Change the values of the primary and secondary
*			DC resistance.
*
* These parameters are underlined.
*
.SUBCKT TRANSF 1 2 3 4
*       ------
* 
LPRIM    5    2    200UH
*                  -----
*
RPS      1    5    5.0
*                  ---
*
LSEC     6    4    200UH
*                  ----
*
RSS      3    6    .001
*                  ----
*
KPS      LPRIM LSEC  .999
*                    ----
.ENDS


.END
